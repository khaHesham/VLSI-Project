
// 	Tue Jan  3 11:09:32 2023
//	vlsi
//	localhost.localdomain

module datapath__0_16 (p_0, adder, p_1);

output [63:0] p_1;
input [63:0] adder;
input [63:0] p_0;
wire n_0;
wire n_367;
wire n_1;
wire n_366;
wire n_365;
wire n_2;
wire n_370;
wire n_364;
wire n_3;
wire n_371;
wire n_376;
wire n_373;
wire n_362;
wire n_10;
wire n_9;
wire n_6;
wire n_7;
wire n_4;
wire n_359;
wire n_350;
wire n_11;
wire n_5;
wire n_360;
wire n_354;
wire n_8;
wire n_357;
wire n_355;
wire n_361;
wire n_352;
wire n_348;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_12;
wire n_345;
wire n_336;
wire n_19;
wire n_13;
wire n_346;
wire n_340;
wire n_16;
wire n_343;
wire n_341;
wire n_347;
wire n_338;
wire n_334;
wire n_26;
wire n_25;
wire n_22;
wire n_23;
wire n_20;
wire n_331;
wire n_322;
wire n_27;
wire n_21;
wire n_332;
wire n_326;
wire n_24;
wire n_329;
wire n_327;
wire n_333;
wire n_324;
wire n_320;
wire n_34;
wire n_33;
wire n_30;
wire n_31;
wire n_28;
wire n_286;
wire n_276;
wire n_35;
wire n_29;
wire n_285;
wire n_288;
wire n_278;
wire n_32;
wire n_287;
wire n_283;
wire n_280;
wire n_290;
wire n_63;
wire n_42;
wire n_41;
wire n_38;
wire n_39;
wire n_36;
wire n_314;
wire n_258;
wire n_43;
wire n_37;
wire n_313;
wire n_316;
wire n_260;
wire n_40;
wire n_315;
wire n_319;
wire n_262;
wire n_318;
wire n_61;
wire n_50;
wire n_49;
wire n_46;
wire n_47;
wire n_44;
wire n_297;
wire n_270;
wire n_51;
wire n_45;
wire n_296;
wire n_299;
wire n_272;
wire n_48;
wire n_298;
wire n_294;
wire n_274;
wire n_301;
wire n_59;
wire n_58;
wire n_57;
wire n_54;
wire n_55;
wire n_52;
wire n_306;
wire n_264;
wire n_65;
wire n_53;
wire n_305;
wire n_308;
wire n_267;
wire n_56;
wire n_307;
wire n_303;
wire n_268;
wire n_60;
wire n_269;
wire n_293;
wire n_62;
wire n_257;
wire n_311;
wire n_64;
wire n_275;
wire n_282;
wire n_309;
wire n_377;
wire n_374;
wire n_255;
wire n_72;
wire n_71;
wire n_68;
wire n_69;
wire n_66;
wire n_224;
wire n_214;
wire n_73;
wire n_67;
wire n_223;
wire n_226;
wire n_216;
wire n_70;
wire n_225;
wire n_221;
wire n_218;
wire n_228;
wire n_101;
wire n_80;
wire n_79;
wire n_76;
wire n_77;
wire n_74;
wire n_249;
wire n_207;
wire n_81;
wire n_75;
wire n_248;
wire n_251;
wire n_209;
wire n_78;
wire n_250;
wire n_254;
wire n_211;
wire n_253;
wire n_99;
wire n_88;
wire n_87;
wire n_84;
wire n_85;
wire n_82;
wire n_235;
wire n_193;
wire n_89;
wire n_83;
wire n_234;
wire n_237;
wire n_195;
wire n_86;
wire n_236;
wire n_232;
wire n_197;
wire n_239;
wire n_98;
wire n_97;
wire n_95;
wire n_94;
wire n_91;
wire n_90;
wire n_203;
wire n_243;
wire n_200;
wire n_103;
wire n_92;
wire n_93;
wire n_242;
wire n_201;
wire n_96;
wire n_244;
wire n_204;
wire n_205;
wire n_192;
wire n_231;
wire n_100;
wire n_206;
wire n_246;
wire n_102;
wire n_213;
wire n_220;
wire n_245;
wire n_190;
wire n_110;
wire n_109;
wire n_106;
wire n_107;
wire n_104;
wire n_187;
wire n_178;
wire n_111;
wire n_105;
wire n_188;
wire n_182;
wire n_108;
wire n_185;
wire n_183;
wire n_189;
wire n_180;
wire n_176;
wire n_118;
wire n_117;
wire n_114;
wire n_115;
wire n_112;
wire n_165;
wire n_155;
wire n_119;
wire n_113;
wire n_164;
wire n_167;
wire n_157;
wire n_116;
wire n_166;
wire n_162;
wire n_159;
wire n_169;
wire n_128;
wire n_127;
wire n_125;
wire n_124;
wire n_121;
wire n_120;
wire n_150;
wire n_173;
wire n_146;
wire n_129;
wire n_122;
wire n_123;
wire n_172;
wire n_147;
wire n_126;
wire n_174;
wire n_151;
wire n_152;
wire n_154;
wire n_161;
wire n_175;
wire n_144;
wire n_143;
wire n_141;
wire n_136;
wire n_142;
wire n_137;
wire n_131;
wire n_130;
wire n_138;
wire n_140;
wire n_133;
wire n_132;
wire n_134;
wire n_135;
wire n_139;
wire n_372;
wire n_148;
wire n_145;
wire n_153;
wire n_160;
wire n_378;
wire n_375;
wire n_149;
wire n_171;
wire n_170;
wire n_156;
wire n_168;
wire n_163;
wire n_158;
wire n_177;
wire n_181;
wire n_184;
wire n_179;
wire n_186;
wire n_212;
wire n_191;
wire n_219;
wire n_198;
wire n_240;
wire n_230;
wire n_194;
wire n_238;
wire n_233;
wire n_196;
wire n_199;
wire n_202;
wire n_241;
wire n_208;
wire n_252;
wire n_247;
wire n_210;
wire n_229;
wire n_215;
wire n_227;
wire n_222;
wire n_217;
wire n_263;
wire n_256;
wire n_281;
wire n_291;
wire n_292;
wire n_302;
wire n_259;
wire n_317;
wire n_312;
wire n_261;
wire n_304;
wire n_266;
wire n_310;
wire n_265;
wire n_271;
wire n_300;
wire n_295;
wire n_273;
wire n_277;
wire n_289;
wire n_284;
wire n_279;
wire n_321;
wire n_325;
wire n_328;
wire n_323;
wire n_330;
wire n_335;
wire n_339;
wire n_342;
wire n_337;
wire n_344;
wire n_349;
wire n_353;
wire n_356;
wire n_351;
wire n_358;
wire n_363;
wire n_369;
wire n_368;


INV_X1 i_442 (.ZN (n_378), .A (p_0[59]));
INV_X1 i_441 (.ZN (n_377), .A (p_0[31]));
INV_X1 i_440 (.ZN (n_376), .A (p_0[3]));
INV_X1 i_439 (.ZN (n_375), .A (adder[59]));
INV_X1 i_438 (.ZN (n_374), .A (adder[31]));
INV_X1 i_437 (.ZN (n_373), .A (adder[3]));
NOR2_X1 i_436 (.ZN (n_372), .A1 (p_0[60]), .A2 (adder[60]));
NAND2_X1 i_435 (.ZN (n_371), .A1 (n_376), .A2 (n_373));
NAND2_X1 i_434 (.ZN (n_370), .A1 (p_0[2]), .A2 (adder[2]));
INV_X1 i_433 (.ZN (n_369), .A (n_370));
NOR2_X1 i_432 (.ZN (n_368), .A1 (p_0[1]), .A2 (adder[1]));
NAND2_X1 i_431 (.ZN (n_367), .A1 (p_0[0]), .A2 (adder[0]));
NAND2_X1 i_430 (.ZN (n_366), .A1 (p_0[1]), .A2 (adder[1]));
AOI21_X1 i_429 (.ZN (n_365), .A (n_368), .B1 (n_367), .B2 (n_366));
OAI22_X1 i_428 (.ZN (n_364), .A1 (p_0[2]), .A2 (adder[2]), .B1 (n_369), .B2 (n_365));
OAI21_X1 i_427 (.ZN (n_363), .A (n_364), .B1 (n_376), .B2 (n_373));
NAND2_X1 i_426 (.ZN (n_362), .A1 (n_371), .A2 (n_363));
NOR2_X1 i_425 (.ZN (n_361), .A1 (p_0[7]), .A2 (adder[7]));
NOR2_X1 i_424 (.ZN (n_360), .A1 (p_0[5]), .A2 (adder[5]));
NOR2_X1 i_423 (.ZN (n_359), .A1 (p_0[6]), .A2 (adder[6]));
OR3_X1 i_422 (.ZN (n_358), .A1 (n_361), .A2 (n_359), .A3 (n_360));
NOR2_X1 i_421 (.ZN (n_357), .A1 (p_0[4]), .A2 (adder[4]));
NOR3_X1 i_420 (.ZN (n_356), .A1 (n_358), .A2 (n_357), .A3 (n_362));
NAND2_X1 i_419 (.ZN (n_355), .A1 (p_0[4]), .A2 (adder[4]));
NAND2_X1 i_418 (.ZN (n_354), .A1 (p_0[5]), .A2 (adder[5]));
AOI21_X1 i_417 (.ZN (n_353), .A (n_358), .B1 (n_355), .B2 (n_354));
AND2_X1 i_416 (.ZN (n_352), .A1 (p_0[7]), .A2 (adder[7]));
NAND2_X1 i_415 (.ZN (n_351), .A1 (p_0[6]), .A2 (adder[6]));
INV_X1 i_414 (.ZN (n_350), .A (n_351));
NOR2_X1 i_413 (.ZN (n_349), .A1 (n_361), .A2 (n_351));
NOR4_X4 i_412 (.ZN (n_348), .A1 (n_352), .A2 (n_349), .A3 (n_353), .A4 (n_356));
NOR2_X1 i_411 (.ZN (n_347), .A1 (p_0[11]), .A2 (adder[11]));
NOR2_X1 i_410 (.ZN (n_346), .A1 (p_0[9]), .A2 (adder[9]));
NOR2_X1 i_409 (.ZN (n_345), .A1 (p_0[10]), .A2 (adder[10]));
OR3_X1 i_408 (.ZN (n_344), .A1 (n_347), .A2 (n_345), .A3 (n_346));
NOR2_X1 i_407 (.ZN (n_343), .A1 (p_0[8]), .A2 (adder[8]));
NOR3_X1 i_406 (.ZN (n_342), .A1 (n_344), .A2 (n_343), .A3 (n_348));
NAND2_X1 i_405 (.ZN (n_341), .A1 (p_0[8]), .A2 (adder[8]));
NAND2_X1 i_404 (.ZN (n_340), .A1 (p_0[9]), .A2 (adder[9]));
AOI21_X1 i_403 (.ZN (n_339), .A (n_344), .B1 (n_341), .B2 (n_340));
AND2_X1 i_402 (.ZN (n_338), .A1 (p_0[11]), .A2 (adder[11]));
NAND2_X1 i_401 (.ZN (n_337), .A1 (p_0[10]), .A2 (adder[10]));
INV_X1 i_400 (.ZN (n_336), .A (n_337));
NOR2_X1 i_399 (.ZN (n_335), .A1 (n_347), .A2 (n_337));
NOR4_X2 i_398 (.ZN (n_334), .A1 (n_338), .A2 (n_335), .A3 (n_339), .A4 (n_342));
NOR2_X1 i_397 (.ZN (n_333), .A1 (p_0[15]), .A2 (adder[15]));
NOR2_X1 i_396 (.ZN (n_332), .A1 (p_0[13]), .A2 (adder[13]));
NOR2_X1 i_395 (.ZN (n_331), .A1 (p_0[14]), .A2 (adder[14]));
OR3_X1 i_394 (.ZN (n_330), .A1 (n_333), .A2 (n_331), .A3 (n_332));
NOR2_X1 i_393 (.ZN (n_329), .A1 (p_0[12]), .A2 (adder[12]));
NOR3_X1 i_392 (.ZN (n_328), .A1 (n_330), .A2 (n_329), .A3 (n_334));
NAND2_X1 i_391 (.ZN (n_327), .A1 (p_0[12]), .A2 (adder[12]));
NAND2_X1 i_390 (.ZN (n_326), .A1 (p_0[13]), .A2 (adder[13]));
AOI21_X1 i_389 (.ZN (n_325), .A (n_330), .B1 (n_327), .B2 (n_326));
AND2_X1 i_388 (.ZN (n_324), .A1 (p_0[15]), .A2 (adder[15]));
NAND2_X1 i_387 (.ZN (n_323), .A1 (p_0[14]), .A2 (adder[14]));
INV_X1 i_386 (.ZN (n_322), .A (n_323));
NOR2_X1 i_385 (.ZN (n_321), .A1 (n_333), .A2 (n_323));
NOR4_X4 i_384 (.ZN (n_320), .A1 (n_324), .A2 (n_321), .A3 (n_325), .A4 (n_328));
NOR2_X1 i_383 (.ZN (n_319), .A1 (p_0[20]), .A2 (adder[20]));
NOR2_X1 i_382 (.ZN (n_318), .A1 (p_0[23]), .A2 (adder[23]));
INV_X1 i_381 (.ZN (n_317), .A (n_318));
NOR2_X1 i_380 (.ZN (n_316), .A1 (p_0[21]), .A2 (adder[21]));
INV_X1 i_379 (.ZN (n_315), .A (n_316));
NOR2_X1 i_378 (.ZN (n_314), .A1 (p_0[22]), .A2 (adder[22]));
INV_X1 i_377 (.ZN (n_313), .A (n_314));
NAND3_X1 i_376 (.ZN (n_312), .A1 (n_317), .A2 (n_313), .A3 (n_315));
OR2_X1 i_375 (.ZN (n_311), .A1 (n_319), .A2 (n_312));
NOR2_X1 i_374 (.ZN (n_310), .A1 (p_0[31]), .A2 (adder[31]));
INV_X1 i_373 (.ZN (n_309), .A (n_310));
NOR2_X1 i_372 (.ZN (n_308), .A1 (p_0[29]), .A2 (adder[29]));
INV_X1 i_371 (.ZN (n_307), .A (n_308));
NOR2_X1 i_370 (.ZN (n_306), .A1 (p_0[30]), .A2 (adder[30]));
INV_X1 i_369 (.ZN (n_305), .A (n_306));
NAND3_X1 i_368 (.ZN (n_304), .A1 (n_309), .A2 (n_305), .A3 (n_307));
NOR2_X1 i_367 (.ZN (n_303), .A1 (p_0[28]), .A2 (adder[28]));
OR2_X1 i_366 (.ZN (n_302), .A1 (n_304), .A2 (n_303));
NOR2_X1 i_365 (.ZN (n_301), .A1 (p_0[27]), .A2 (adder[27]));
INV_X1 i_364 (.ZN (n_300), .A (n_301));
NOR2_X1 i_363 (.ZN (n_299), .A1 (p_0[25]), .A2 (adder[25]));
INV_X1 i_362 (.ZN (n_298), .A (n_299));
NOR2_X1 i_361 (.ZN (n_297), .A1 (p_0[26]), .A2 (adder[26]));
INV_X1 i_360 (.ZN (n_296), .A (n_297));
NAND3_X1 i_359 (.ZN (n_295), .A1 (n_300), .A2 (n_296), .A3 (n_298));
NOR2_X1 i_358 (.ZN (n_294), .A1 (p_0[24]), .A2 (adder[24]));
OR2_X1 i_357 (.ZN (n_293), .A1 (n_295), .A2 (n_294));
OR2_X1 i_356 (.ZN (n_292), .A1 (n_302), .A2 (n_293));
OR2_X1 i_355 (.ZN (n_291), .A1 (n_311), .A2 (n_292));
NOR2_X1 i_354 (.ZN (n_290), .A1 (p_0[19]), .A2 (adder[19]));
INV_X1 i_353 (.ZN (n_289), .A (n_290));
NOR2_X1 i_352 (.ZN (n_288), .A1 (p_0[17]), .A2 (adder[17]));
INV_X1 i_351 (.ZN (n_287), .A (n_288));
NOR2_X1 i_350 (.ZN (n_286), .A1 (p_0[18]), .A2 (adder[18]));
INV_X1 i_349 (.ZN (n_285), .A (n_286));
NAND3_X1 i_348 (.ZN (n_284), .A1 (n_289), .A2 (n_285), .A3 (n_287));
NOR2_X1 i_347 (.ZN (n_283), .A1 (p_0[16]), .A2 (adder[16]));
OR2_X1 i_346 (.ZN (n_282), .A1 (n_284), .A2 (n_283));
NOR3_X1 i_345 (.ZN (n_281), .A1 (n_291), .A2 (n_282), .A3 (n_320));
NAND2_X1 i_344 (.ZN (n_280), .A1 (p_0[16]), .A2 (adder[16]));
NAND2_X1 i_343 (.ZN (n_279), .A1 (p_0[17]), .A2 (adder[17]));
INV_X1 i_342 (.ZN (n_278), .A (n_279));
AOI21_X1 i_341 (.ZN (n_277), .A (n_284), .B1 (n_280), .B2 (n_279));
AND2_X1 i_340 (.ZN (n_276), .A1 (p_0[18]), .A2 (adder[18]));
AOI221_X1 i_339 (.ZN (n_275), .A (n_277), .B1 (p_0[19]), .B2 (adder[19]), .C1 (n_289), .C2 (n_276));
NAND2_X1 i_338 (.ZN (n_274), .A1 (p_0[24]), .A2 (adder[24]));
NAND2_X1 i_337 (.ZN (n_273), .A1 (p_0[25]), .A2 (adder[25]));
INV_X1 i_336 (.ZN (n_272), .A (n_273));
AOI21_X1 i_335 (.ZN (n_271), .A (n_295), .B1 (n_274), .B2 (n_273));
AND2_X1 i_334 (.ZN (n_270), .A1 (p_0[26]), .A2 (adder[26]));
AOI221_X1 i_333 (.ZN (n_269), .A (n_271), .B1 (p_0[27]), .B2 (adder[27]), .C1 (n_300), .C2 (n_270));
NAND2_X1 i_332 (.ZN (n_268), .A1 (p_0[28]), .A2 (adder[28]));
AND2_X1 i_331 (.ZN (n_267), .A1 (p_0[29]), .A2 (adder[29]));
AOI21_X1 i_330 (.ZN (n_266), .A (n_267), .B1 (p_0[28]), .B2 (adder[28]));
NAND2_X1 i_329 (.ZN (n_265), .A1 (p_0[30]), .A2 (adder[30]));
INV_X1 i_328 (.ZN (n_264), .A (n_265));
OAI222_X1 i_327 (.ZN (n_263), .A1 (n_304), .A2 (n_266), .B1 (n_310), .B2 (n_265), .C1 (n_377), .C2 (n_374));
NAND2_X1 i_326 (.ZN (n_262), .A1 (p_0[20]), .A2 (adder[20]));
NAND2_X1 i_325 (.ZN (n_261), .A1 (p_0[21]), .A2 (adder[21]));
INV_X1 i_324 (.ZN (n_260), .A (n_261));
AOI21_X1 i_323 (.ZN (n_259), .A (n_312), .B1 (n_262), .B2 (n_261));
AND2_X1 i_322 (.ZN (n_258), .A1 (p_0[22]), .A2 (adder[22]));
AOI221_X1 i_321 (.ZN (n_257), .A (n_259), .B1 (p_0[23]), .B2 (adder[23]), .C1 (n_317), .C2 (n_258));
OAI222_X1 i_320 (.ZN (n_256), .A1 (n_291), .A2 (n_275), .B1 (n_292), .B2 (n_257), .C1 (n_302), .C2 (n_269));
NOR3_X4 i_319 (.ZN (n_255), .A1 (n_263), .A2 (n_256), .A3 (n_281));
NOR2_X1 i_318 (.ZN (n_254), .A1 (p_0[36]), .A2 (adder[36]));
NOR2_X1 i_317 (.ZN (n_253), .A1 (p_0[39]), .A2 (adder[39]));
INV_X1 i_316 (.ZN (n_252), .A (n_253));
NOR2_X1 i_315 (.ZN (n_251), .A1 (p_0[37]), .A2 (adder[37]));
INV_X1 i_314 (.ZN (n_250), .A (n_251));
NOR2_X1 i_313 (.ZN (n_249), .A1 (p_0[38]), .A2 (adder[38]));
INV_X1 i_312 (.ZN (n_248), .A (n_249));
NAND3_X1 i_311 (.ZN (n_247), .A1 (n_252), .A2 (n_248), .A3 (n_250));
OR2_X1 i_310 (.ZN (n_246), .A1 (n_254), .A2 (n_247));
NOR2_X1 i_309 (.ZN (n_245), .A1 (p_0[47]), .A2 (adder[47]));
NOR2_X1 i_308 (.ZN (n_244), .A1 (p_0[45]), .A2 (adder[45]));
NOR2_X1 i_307 (.ZN (n_243), .A1 (p_0[46]), .A2 (adder[46]));
NOR2_X1 i_306 (.ZN (n_242), .A1 (n_244), .A2 (n_243));
NOR3_X1 i_305 (.ZN (n_241), .A1 (n_245), .A2 (n_243), .A3 (n_244));
OAI21_X1 i_304 (.ZN (n_240), .A (n_241), .B1 (p_0[44]), .B2 (adder[44]));
NOR2_X1 i_303 (.ZN (n_239), .A1 (p_0[43]), .A2 (adder[43]));
INV_X1 i_302 (.ZN (n_238), .A (n_239));
NOR2_X1 i_301 (.ZN (n_237), .A1 (p_0[41]), .A2 (adder[41]));
INV_X1 i_300 (.ZN (n_236), .A (n_237));
NOR2_X1 i_299 (.ZN (n_235), .A1 (p_0[42]), .A2 (adder[42]));
INV_X1 i_298 (.ZN (n_234), .A (n_235));
NAND3_X1 i_297 (.ZN (n_233), .A1 (n_238), .A2 (n_234), .A3 (n_236));
NOR2_X1 i_296 (.ZN (n_232), .A1 (p_0[40]), .A2 (adder[40]));
OR2_X1 i_295 (.ZN (n_231), .A1 (n_233), .A2 (n_232));
OR2_X1 i_294 (.ZN (n_230), .A1 (n_240), .A2 (n_231));
OR2_X1 i_293 (.ZN (n_229), .A1 (n_246), .A2 (n_230));
NOR2_X1 i_292 (.ZN (n_228), .A1 (p_0[35]), .A2 (adder[35]));
INV_X1 i_291 (.ZN (n_227), .A (n_228));
NOR2_X1 i_290 (.ZN (n_226), .A1 (p_0[33]), .A2 (adder[33]));
INV_X1 i_289 (.ZN (n_225), .A (n_226));
NOR2_X1 i_288 (.ZN (n_224), .A1 (p_0[34]), .A2 (adder[34]));
INV_X1 i_287 (.ZN (n_223), .A (n_224));
NAND3_X1 i_286 (.ZN (n_222), .A1 (n_227), .A2 (n_223), .A3 (n_225));
NOR2_X1 i_285 (.ZN (n_221), .A1 (p_0[32]), .A2 (adder[32]));
OR2_X1 i_284 (.ZN (n_220), .A1 (n_222), .A2 (n_221));
NOR3_X1 i_283 (.ZN (n_219), .A1 (n_229), .A2 (n_220), .A3 (n_255));
NAND2_X1 i_282 (.ZN (n_218), .A1 (p_0[32]), .A2 (adder[32]));
NAND2_X1 i_281 (.ZN (n_217), .A1 (p_0[33]), .A2 (adder[33]));
INV_X1 i_280 (.ZN (n_216), .A (n_217));
AOI21_X1 i_279 (.ZN (n_215), .A (n_222), .B1 (n_218), .B2 (n_217));
AND2_X1 i_278 (.ZN (n_214), .A1 (p_0[34]), .A2 (adder[34]));
AOI221_X1 i_277 (.ZN (n_213), .A (n_215), .B1 (p_0[35]), .B2 (adder[35]), .C1 (n_227), .C2 (n_214));
NOR2_X1 i_276 (.ZN (n_212), .A1 (n_229), .A2 (n_213));
NAND2_X1 i_275 (.ZN (n_211), .A1 (p_0[36]), .A2 (adder[36]));
NAND2_X1 i_274 (.ZN (n_210), .A1 (p_0[37]), .A2 (adder[37]));
INV_X1 i_273 (.ZN (n_209), .A (n_210));
AOI21_X1 i_272 (.ZN (n_208), .A (n_247), .B1 (n_211), .B2 (n_210));
AND2_X1 i_271 (.ZN (n_207), .A1 (p_0[38]), .A2 (adder[38]));
AOI221_X1 i_270 (.ZN (n_206), .A (n_208), .B1 (p_0[39]), .B2 (adder[39]), .C1 (n_252), .C2 (n_207));
NAND2_X1 i_269 (.ZN (n_205), .A1 (p_0[44]), .A2 (adder[44]));
INV_X1 i_268 (.ZN (n_204), .A (n_205));
AND2_X1 i_267 (.ZN (n_203), .A1 (p_0[45]), .A2 (adder[45]));
OAI21_X1 i_266 (.ZN (n_202), .A (n_241), .B1 (n_204), .B2 (n_203));
NAND2_X1 i_265 (.ZN (n_201), .A1 (p_0[46]), .A2 (adder[46]));
INV_X1 i_264 (.ZN (n_200), .A (n_201));
OAI21_X1 i_263 (.ZN (n_199), .A (n_202), .B1 (n_245), .B2 (n_201));
AOI21_X1 i_262 (.ZN (n_198), .A (n_199), .B1 (p_0[47]), .B2 (adder[47]));
NAND2_X1 i_261 (.ZN (n_197), .A1 (p_0[40]), .A2 (adder[40]));
NAND2_X1 i_260 (.ZN (n_196), .A1 (p_0[41]), .A2 (adder[41]));
INV_X1 i_259 (.ZN (n_195), .A (n_196));
AOI21_X1 i_258 (.ZN (n_194), .A (n_233), .B1 (n_197), .B2 (n_196));
AND2_X1 i_257 (.ZN (n_193), .A1 (p_0[42]), .A2 (adder[42]));
AOI221_X1 i_256 (.ZN (n_192), .A (n_194), .B1 (p_0[43]), .B2 (adder[43]), .C1 (n_238), .C2 (n_193));
OAI221_X1 i_255 (.ZN (n_191), .A (n_198), .B1 (n_240), .B2 (n_192), .C1 (n_230), .C2 (n_206));
NOR3_X1 i_254 (.ZN (n_190), .A1 (n_212), .A2 (n_191), .A3 (n_219));
NOR2_X1 i_253 (.ZN (n_189), .A1 (p_0[51]), .A2 (adder[51]));
NOR2_X1 i_252 (.ZN (n_188), .A1 (p_0[49]), .A2 (adder[49]));
NOR2_X1 i_251 (.ZN (n_187), .A1 (p_0[50]), .A2 (adder[50]));
OR3_X1 i_250 (.ZN (n_186), .A1 (n_189), .A2 (n_187), .A3 (n_188));
NOR2_X1 i_249 (.ZN (n_185), .A1 (p_0[48]), .A2 (adder[48]));
NOR3_X1 i_248 (.ZN (n_184), .A1 (n_186), .A2 (n_185), .A3 (n_190));
NAND2_X1 i_247 (.ZN (n_183), .A1 (p_0[48]), .A2 (adder[48]));
NAND2_X1 i_246 (.ZN (n_182), .A1 (p_0[49]), .A2 (adder[49]));
AOI21_X1 i_245 (.ZN (n_181), .A (n_186), .B1 (n_183), .B2 (n_182));
AND2_X1 i_244 (.ZN (n_180), .A1 (p_0[51]), .A2 (adder[51]));
NAND2_X1 i_243 (.ZN (n_179), .A1 (p_0[50]), .A2 (adder[50]));
INV_X1 i_242 (.ZN (n_178), .A (n_179));
NOR2_X1 i_241 (.ZN (n_177), .A1 (n_189), .A2 (n_179));
NOR4_X4 i_240 (.ZN (n_176), .A1 (n_180), .A2 (n_177), .A3 (n_181), .A4 (n_184));
NOR2_X1 i_239 (.ZN (n_175), .A1 (p_0[59]), .A2 (adder[59]));
NOR2_X1 i_238 (.ZN (n_174), .A1 (p_0[57]), .A2 (adder[57]));
NOR2_X1 i_237 (.ZN (n_173), .A1 (p_0[58]), .A2 (adder[58]));
NOR2_X1 i_236 (.ZN (n_172), .A1 (n_174), .A2 (n_173));
NOR3_X1 i_235 (.ZN (n_171), .A1 (n_175), .A2 (n_173), .A3 (n_174));
OAI21_X1 i_234 (.ZN (n_170), .A (n_171), .B1 (p_0[56]), .B2 (adder[56]));
NOR2_X1 i_233 (.ZN (n_169), .A1 (p_0[55]), .A2 (adder[55]));
INV_X1 i_232 (.ZN (n_168), .A (n_169));
NOR2_X1 i_231 (.ZN (n_167), .A1 (p_0[53]), .A2 (adder[53]));
INV_X1 i_230 (.ZN (n_166), .A (n_167));
NOR2_X1 i_229 (.ZN (n_165), .A1 (p_0[54]), .A2 (adder[54]));
INV_X1 i_228 (.ZN (n_164), .A (n_165));
NAND3_X1 i_227 (.ZN (n_163), .A1 (n_168), .A2 (n_164), .A3 (n_166));
NOR2_X1 i_226 (.ZN (n_162), .A1 (p_0[52]), .A2 (adder[52]));
OR2_X1 i_225 (.ZN (n_161), .A1 (n_163), .A2 (n_162));
NOR3_X1 i_224 (.ZN (n_160), .A1 (n_170), .A2 (n_161), .A3 (n_176));
NAND2_X1 i_223 (.ZN (n_159), .A1 (p_0[52]), .A2 (adder[52]));
NAND2_X1 i_222 (.ZN (n_158), .A1 (p_0[53]), .A2 (adder[53]));
INV_X1 i_221 (.ZN (n_157), .A (n_158));
AOI21_X1 i_220 (.ZN (n_156), .A (n_163), .B1 (n_159), .B2 (n_158));
AND2_X1 i_219 (.ZN (n_155), .A1 (p_0[54]), .A2 (adder[54]));
AOI221_X1 i_218 (.ZN (n_154), .A (n_156), .B1 (p_0[55]), .B2 (adder[55]), .C1 (n_168), .C2 (n_155));
NOR2_X1 i_217 (.ZN (n_153), .A1 (n_170), .A2 (n_154));
NAND2_X1 i_216 (.ZN (n_152), .A1 (p_0[56]), .A2 (adder[56]));
INV_X1 i_215 (.ZN (n_151), .A (n_152));
AND2_X1 i_214 (.ZN (n_150), .A1 (p_0[57]), .A2 (adder[57]));
OAI21_X1 i_213 (.ZN (n_149), .A (n_171), .B1 (n_151), .B2 (n_150));
INV_X1 i_212 (.ZN (n_148), .A (n_149));
NAND2_X1 i_211 (.ZN (n_147), .A1 (p_0[58]), .A2 (adder[58]));
INV_X1 i_210 (.ZN (n_146), .A (n_147));
OAI22_X1 i_209 (.ZN (n_145), .A1 (n_378), .A2 (n_375), .B1 (n_175), .B2 (n_147));
NOR4_X1 i_208 (.ZN (n_144), .A1 (n_148), .A2 (n_145), .A3 (n_153), .A4 (n_160));
AOI21_X1 i_207 (.ZN (n_143), .A (n_372), .B1 (p_0[60]), .B2 (adder[60]));
AOI21_X1 i_206 (.ZN (n_142), .A (n_372), .B1 (n_144), .B2 (n_143));
INV_X1 i_205 (.ZN (n_141), .A (n_142));
NOR2_X1 i_204 (.ZN (n_140), .A1 (p_0[61]), .A2 (adder[62]));
NOR2_X1 i_203 (.ZN (n_139), .A1 (p_0[61]), .A2 (adder[61]));
INV_X1 i_202 (.ZN (n_138), .A (n_139));
AOI21_X1 i_201 (.ZN (n_137), .A (n_139), .B1 (p_0[61]), .B2 (adder[61]));
INV_X1 i_200 (.ZN (n_136), .A (n_137));
NOR2_X1 i_199 (.ZN (n_135), .A1 (n_140), .A2 (n_136));
NOR2_X1 i_198 (.ZN (n_134), .A1 (n_140), .A2 (n_138));
AOI221_X1 i_197 (.ZN (n_133), .A (n_134), .B1 (p_0[61]), .B2 (adder[62]), .C1 (n_141), .C2 (n_135));
XOR2_X1 i_196 (.Z (n_132), .A (adder[63]), .B (adder[62]));
XNOR2_X1 i_195 (.ZN (p_1[63]), .A (n_133), .B (n_132));
AOI21_X1 i_194 (.ZN (n_131), .A (n_140), .B1 (p_0[61]), .B2 (adder[62]));
AOI22_X1 i_193 (.ZN (n_130), .A1 (p_0[61]), .A2 (adder[61]), .B1 (n_142), .B2 (n_138));
XNOR2_X1 i_192 (.ZN (p_1[62]), .A (n_131), .B (n_130));
AOI22_X1 i_191 (.ZN (p_1[61]), .A1 (n_141), .A2 (n_136), .B1 (n_142), .B2 (n_137));
XNOR2_X1 i_190 (.ZN (p_1[60]), .A (n_144), .B (n_143));
AOI21_X1 i_189 (.ZN (n_129), .A (n_175), .B1 (p_0[59]), .B2 (adder[59]));
OAI21_X1 i_188 (.ZN (n_128), .A (n_154), .B1 (n_176), .B2 (n_161));
OAI21_X1 i_187 (.ZN (n_127), .A (n_152), .B1 (p_0[56]), .B2 (adder[56]));
OAI22_X1 i_186 (.ZN (n_126), .A1 (p_0[56]), .A2 (adder[56]), .B1 (n_151), .B2 (n_128));
INV_X1 i_185 (.ZN (n_125), .A (n_126));
NOR2_X1 i_184 (.ZN (n_124), .A1 (n_174), .A2 (n_150));
NAND3_X1 i_183 (.ZN (n_123), .A1 (n_147), .A2 (n_124), .A3 (n_126));
OAI21_X1 i_182 (.ZN (n_122), .A (n_123), .B1 (n_172), .B2 (n_146));
XNOR2_X1 i_181 (.ZN (p_1[59]), .A (n_129), .B (n_122));
NOR2_X1 i_180 (.ZN (n_121), .A1 (n_173), .A2 (n_146));
OAI22_X1 i_179 (.ZN (n_120), .A1 (p_0[57]), .A2 (adder[57]), .B1 (n_150), .B2 (n_125));
XNOR2_X1 i_178 (.ZN (p_1[58]), .A (n_121), .B (n_120));
XOR2_X1 i_177 (.Z (p_1[57]), .A (n_125), .B (n_124));
XNOR2_X1 i_176 (.ZN (p_1[56]), .A (n_128), .B (n_127));
AOI21_X1 i_175 (.ZN (n_119), .A (n_169), .B1 (p_0[55]), .B2 (adder[55]));
OAI21_X1 i_174 (.ZN (n_118), .A (n_159), .B1 (p_0[52]), .B2 (adder[52]));
AOI21_X1 i_173 (.ZN (n_117), .A (n_162), .B1 (n_176), .B2 (n_159));
OAI21_X1 i_172 (.ZN (n_116), .A (n_166), .B1 (n_157), .B2 (n_117));
INV_X1 i_171 (.ZN (n_115), .A (n_116));
NOR2_X1 i_170 (.ZN (n_114), .A1 (n_167), .A2 (n_157));
OAI21_X1 i_169 (.ZN (n_113), .A (n_164), .B1 (n_155), .B2 (n_115));
XNOR2_X1 i_168 (.ZN (p_1[55]), .A (n_119), .B (n_113));
NOR2_X1 i_167 (.ZN (n_112), .A1 (n_165), .A2 (n_155));
XOR2_X1 i_166 (.Z (p_1[54]), .A (n_115), .B (n_112));
XOR2_X1 i_165 (.Z (p_1[53]), .A (n_117), .B (n_114));
XOR2_X1 i_164 (.Z (p_1[52]), .A (n_176), .B (n_118));
NOR2_X1 i_163 (.ZN (n_111), .A1 (n_189), .A2 (n_180));
OAI21_X1 i_162 (.ZN (n_110), .A (n_183), .B1 (p_0[48]), .B2 (adder[48]));
AOI21_X1 i_161 (.ZN (n_109), .A (n_185), .B1 (n_190), .B2 (n_183));
INV_X1 i_160 (.ZN (n_108), .A (n_109));
AOI21_X1 i_159 (.ZN (n_107), .A (n_188), .B1 (n_182), .B2 (n_108));
AOI21_X1 i_158 (.ZN (n_106), .A (n_188), .B1 (p_0[49]), .B2 (adder[49]));
OAI22_X1 i_157 (.ZN (n_105), .A1 (p_0[50]), .A2 (adder[50]), .B1 (n_178), .B2 (n_107));
XNOR2_X1 i_156 (.ZN (p_1[51]), .A (n_111), .B (n_105));
NOR2_X1 i_155 (.ZN (n_104), .A1 (n_187), .A2 (n_178));
XOR2_X1 i_154 (.Z (p_1[50]), .A (n_107), .B (n_104));
XOR2_X1 i_153 (.Z (p_1[49]), .A (n_109), .B (n_106));
XOR2_X1 i_152 (.Z (p_1[48]), .A (n_190), .B (n_110));
AOI21_X1 i_151 (.ZN (n_103), .A (n_245), .B1 (p_0[47]), .B2 (adder[47]));
OAI21_X1 i_150 (.ZN (n_102), .A (n_213), .B1 (n_255), .B2 (n_220));
INV_X1 i_149 (.ZN (n_101), .A (n_102));
OAI21_X1 i_148 (.ZN (n_100), .A (n_206), .B1 (n_246), .B2 (n_101));
INV_X1 i_147 (.ZN (n_99), .A (n_100));
OAI21_X1 i_146 (.ZN (n_98), .A (n_192), .B1 (n_231), .B2 (n_99));
OAI21_X1 i_145 (.ZN (n_97), .A (n_205), .B1 (p_0[44]), .B2 (adder[44]));
OAI22_X1 i_144 (.ZN (n_96), .A1 (p_0[44]), .A2 (adder[44]), .B1 (n_204), .B2 (n_98));
INV_X1 i_143 (.ZN (n_95), .A (n_96));
NOR2_X1 i_142 (.ZN (n_94), .A1 (n_244), .A2 (n_203));
NAND3_X1 i_141 (.ZN (n_93), .A1 (n_201), .A2 (n_94), .A3 (n_96));
OAI21_X1 i_140 (.ZN (n_92), .A (n_93), .B1 (n_242), .B2 (n_200));
XNOR2_X1 i_139 (.ZN (p_1[47]), .A (n_103), .B (n_92));
NOR2_X1 i_138 (.ZN (n_91), .A1 (n_243), .A2 (n_200));
OAI22_X1 i_137 (.ZN (n_90), .A1 (p_0[45]), .A2 (adder[45]), .B1 (n_203), .B2 (n_95));
XNOR2_X1 i_136 (.ZN (p_1[46]), .A (n_91), .B (n_90));
XOR2_X1 i_135 (.Z (p_1[45]), .A (n_95), .B (n_94));
XNOR2_X1 i_134 (.ZN (p_1[44]), .A (n_98), .B (n_97));
AOI21_X1 i_133 (.ZN (n_89), .A (n_239), .B1 (p_0[43]), .B2 (adder[43]));
OAI21_X1 i_132 (.ZN (n_88), .A (n_197), .B1 (p_0[40]), .B2 (adder[40]));
AOI21_X1 i_131 (.ZN (n_87), .A (n_232), .B1 (n_197), .B2 (n_99));
OAI21_X1 i_130 (.ZN (n_86), .A (n_236), .B1 (n_195), .B2 (n_87));
INV_X1 i_129 (.ZN (n_85), .A (n_86));
NOR2_X1 i_128 (.ZN (n_84), .A1 (n_237), .A2 (n_195));
OAI21_X1 i_127 (.ZN (n_83), .A (n_234), .B1 (n_193), .B2 (n_85));
XNOR2_X1 i_126 (.ZN (p_1[43]), .A (n_89), .B (n_83));
NOR2_X1 i_125 (.ZN (n_82), .A1 (n_235), .A2 (n_193));
XOR2_X1 i_124 (.Z (p_1[42]), .A (n_85), .B (n_82));
XOR2_X1 i_123 (.Z (p_1[41]), .A (n_87), .B (n_84));
XOR2_X1 i_122 (.Z (p_1[40]), .A (n_99), .B (n_88));
AOI21_X1 i_121 (.ZN (n_81), .A (n_253), .B1 (p_0[39]), .B2 (adder[39]));
OAI21_X1 i_120 (.ZN (n_80), .A (n_211), .B1 (p_0[36]), .B2 (adder[36]));
AOI21_X1 i_119 (.ZN (n_79), .A (n_254), .B1 (n_211), .B2 (n_101));
OAI21_X1 i_118 (.ZN (n_78), .A (n_250), .B1 (n_209), .B2 (n_79));
INV_X1 i_117 (.ZN (n_77), .A (n_78));
NOR2_X1 i_116 (.ZN (n_76), .A1 (n_251), .A2 (n_209));
OAI21_X1 i_115 (.ZN (n_75), .A (n_248), .B1 (n_207), .B2 (n_77));
XNOR2_X1 i_114 (.ZN (p_1[39]), .A (n_81), .B (n_75));
NOR2_X1 i_113 (.ZN (n_74), .A1 (n_249), .A2 (n_207));
XOR2_X1 i_112 (.Z (p_1[38]), .A (n_77), .B (n_74));
XOR2_X1 i_111 (.Z (p_1[37]), .A (n_79), .B (n_76));
XOR2_X1 i_110 (.Z (p_1[36]), .A (n_101), .B (n_80));
AOI21_X1 i_109 (.ZN (n_73), .A (n_228), .B1 (p_0[35]), .B2 (adder[35]));
OAI21_X1 i_108 (.ZN (n_72), .A (n_218), .B1 (p_0[32]), .B2 (adder[32]));
AOI21_X1 i_107 (.ZN (n_71), .A (n_221), .B1 (n_255), .B2 (n_218));
OAI21_X1 i_106 (.ZN (n_70), .A (n_225), .B1 (n_216), .B2 (n_71));
INV_X1 i_105 (.ZN (n_69), .A (n_70));
NOR2_X1 i_104 (.ZN (n_68), .A1 (n_226), .A2 (n_216));
OAI21_X1 i_103 (.ZN (n_67), .A (n_223), .B1 (n_214), .B2 (n_69));
XNOR2_X1 i_102 (.ZN (p_1[35]), .A (n_73), .B (n_67));
NOR2_X1 i_101 (.ZN (n_66), .A1 (n_224), .A2 (n_214));
XOR2_X1 i_100 (.Z (p_1[34]), .A (n_69), .B (n_66));
XOR2_X1 i_99 (.Z (p_1[33]), .A (n_71), .B (n_68));
XOR2_X1 i_98 (.Z (p_1[32]), .A (n_255), .B (n_72));
OAI21_X1 i_97 (.ZN (n_65), .A (n_309), .B1 (n_377), .B2 (n_374));
OAI21_X1 i_96 (.ZN (n_64), .A (n_275), .B1 (n_320), .B2 (n_282));
INV_X1 i_95 (.ZN (n_63), .A (n_64));
OAI21_X1 i_94 (.ZN (n_62), .A (n_257), .B1 (n_311), .B2 (n_63));
INV_X1 i_93 (.ZN (n_61), .A (n_62));
OAI21_X1 i_92 (.ZN (n_60), .A (n_269), .B1 (n_293), .B2 (n_61));
INV_X1 i_91 (.ZN (n_59), .A (n_60));
OAI21_X1 i_90 (.ZN (n_58), .A (n_268), .B1 (p_0[28]), .B2 (adder[28]));
AOI21_X1 i_89 (.ZN (n_57), .A (n_303), .B1 (n_268), .B2 (n_59));
OAI21_X1 i_88 (.ZN (n_56), .A (n_307), .B1 (n_267), .B2 (n_57));
INV_X1 i_87 (.ZN (n_55), .A (n_56));
NOR2_X1 i_86 (.ZN (n_54), .A1 (n_308), .A2 (n_267));
OAI21_X1 i_85 (.ZN (n_53), .A (n_305), .B1 (n_264), .B2 (n_55));
XOR2_X1 i_84 (.Z (p_1[31]), .A (n_65), .B (n_53));
NOR2_X1 i_83 (.ZN (n_52), .A1 (n_306), .A2 (n_264));
XOR2_X1 i_82 (.Z (p_1[30]), .A (n_55), .B (n_52));
XOR2_X1 i_81 (.Z (p_1[29]), .A (n_57), .B (n_54));
XOR2_X1 i_80 (.Z (p_1[28]), .A (n_59), .B (n_58));
AOI21_X1 i_79 (.ZN (n_51), .A (n_301), .B1 (p_0[27]), .B2 (adder[27]));
OAI21_X1 i_78 (.ZN (n_50), .A (n_274), .B1 (p_0[24]), .B2 (adder[24]));
AOI21_X1 i_77 (.ZN (n_49), .A (n_294), .B1 (n_274), .B2 (n_61));
OAI21_X1 i_76 (.ZN (n_48), .A (n_298), .B1 (n_272), .B2 (n_49));
INV_X1 i_75 (.ZN (n_47), .A (n_48));
NOR2_X1 i_74 (.ZN (n_46), .A1 (n_299), .A2 (n_272));
OAI21_X1 i_73 (.ZN (n_45), .A (n_296), .B1 (n_270), .B2 (n_47));
XNOR2_X1 i_72 (.ZN (p_1[27]), .A (n_51), .B (n_45));
NOR2_X1 i_71 (.ZN (n_44), .A1 (n_297), .A2 (n_270));
XOR2_X1 i_70 (.Z (p_1[26]), .A (n_47), .B (n_44));
XOR2_X1 i_69 (.Z (p_1[25]), .A (n_49), .B (n_46));
XOR2_X1 i_68 (.Z (p_1[24]), .A (n_61), .B (n_50));
AOI21_X1 i_67 (.ZN (n_43), .A (n_318), .B1 (p_0[23]), .B2 (adder[23]));
OAI21_X1 i_66 (.ZN (n_42), .A (n_262), .B1 (p_0[20]), .B2 (adder[20]));
AOI21_X1 i_65 (.ZN (n_41), .A (n_319), .B1 (n_262), .B2 (n_63));
OAI21_X1 i_64 (.ZN (n_40), .A (n_315), .B1 (n_260), .B2 (n_41));
INV_X1 i_63 (.ZN (n_39), .A (n_40));
NOR2_X1 i_62 (.ZN (n_38), .A1 (n_316), .A2 (n_260));
OAI21_X1 i_61 (.ZN (n_37), .A (n_313), .B1 (n_258), .B2 (n_39));
XNOR2_X1 i_60 (.ZN (p_1[23]), .A (n_43), .B (n_37));
NOR2_X1 i_59 (.ZN (n_36), .A1 (n_314), .A2 (n_258));
XOR2_X1 i_58 (.Z (p_1[22]), .A (n_39), .B (n_36));
XOR2_X1 i_57 (.Z (p_1[21]), .A (n_41), .B (n_38));
XOR2_X1 i_56 (.Z (p_1[20]), .A (n_63), .B (n_42));
AOI21_X1 i_55 (.ZN (n_35), .A (n_290), .B1 (p_0[19]), .B2 (adder[19]));
OAI21_X1 i_54 (.ZN (n_34), .A (n_280), .B1 (p_0[16]), .B2 (adder[16]));
AOI21_X1 i_53 (.ZN (n_33), .A (n_283), .B1 (n_320), .B2 (n_280));
OAI21_X1 i_52 (.ZN (n_32), .A (n_287), .B1 (n_278), .B2 (n_33));
INV_X1 i_51 (.ZN (n_31), .A (n_32));
NOR2_X1 i_50 (.ZN (n_30), .A1 (n_288), .A2 (n_278));
OAI21_X1 i_49 (.ZN (n_29), .A (n_285), .B1 (n_276), .B2 (n_31));
XNOR2_X1 i_48 (.ZN (p_1[19]), .A (n_35), .B (n_29));
NOR2_X1 i_47 (.ZN (n_28), .A1 (n_286), .A2 (n_276));
XOR2_X1 i_46 (.Z (p_1[18]), .A (n_31), .B (n_28));
XOR2_X1 i_45 (.Z (p_1[17]), .A (n_33), .B (n_30));
XOR2_X1 i_44 (.Z (p_1[16]), .A (n_320), .B (n_34));
NOR2_X1 i_43 (.ZN (n_27), .A1 (n_333), .A2 (n_324));
OAI21_X1 i_42 (.ZN (n_26), .A (n_327), .B1 (p_0[12]), .B2 (adder[12]));
AOI21_X1 i_41 (.ZN (n_25), .A (n_329), .B1 (n_334), .B2 (n_327));
INV_X1 i_40 (.ZN (n_24), .A (n_25));
AOI21_X1 i_39 (.ZN (n_23), .A (n_332), .B1 (n_326), .B2 (n_24));
AOI21_X1 i_38 (.ZN (n_22), .A (n_332), .B1 (p_0[13]), .B2 (adder[13]));
OAI22_X1 i_37 (.ZN (n_21), .A1 (p_0[14]), .A2 (adder[14]), .B1 (n_322), .B2 (n_23));
XNOR2_X1 i_36 (.ZN (p_1[15]), .A (n_27), .B (n_21));
NOR2_X1 i_35 (.ZN (n_20), .A1 (n_331), .A2 (n_322));
XOR2_X1 i_34 (.Z (p_1[14]), .A (n_23), .B (n_20));
XOR2_X1 i_33 (.Z (p_1[13]), .A (n_25), .B (n_22));
XOR2_X1 i_32 (.Z (p_1[12]), .A (n_334), .B (n_26));
NOR2_X1 i_31 (.ZN (n_19), .A1 (n_347), .A2 (n_338));
AOI21_X1 i_30 (.ZN (n_18), .A (n_343), .B1 (p_0[8]), .B2 (adder[8]));
AOI21_X1 i_29 (.ZN (n_17), .A (n_343), .B1 (n_348), .B2 (n_341));
INV_X1 i_28 (.ZN (n_16), .A (n_17));
AOI21_X1 i_27 (.ZN (n_15), .A (n_346), .B1 (n_340), .B2 (n_16));
AOI21_X1 i_26 (.ZN (n_14), .A (n_346), .B1 (p_0[9]), .B2 (adder[9]));
OAI22_X1 i_25 (.ZN (n_13), .A1 (p_0[10]), .A2 (adder[10]), .B1 (n_336), .B2 (n_15));
XNOR2_X1 i_24 (.ZN (p_1[11]), .A (n_19), .B (n_13));
NOR2_X1 i_23 (.ZN (n_12), .A1 (n_345), .A2 (n_336));
XOR2_X1 i_22 (.Z (p_1[10]), .A (n_15), .B (n_12));
XOR2_X1 i_21 (.Z (p_1[9]), .A (n_17), .B (n_14));
XNOR2_X1 i_20 (.ZN (p_1[8]), .A (n_348), .B (n_18));
NOR2_X1 i_19 (.ZN (n_11), .A1 (n_361), .A2 (n_352));
OAI21_X1 i_18 (.ZN (n_10), .A (n_355), .B1 (p_0[4]), .B2 (adder[4]));
AOI21_X1 i_17 (.ZN (n_9), .A (n_357), .B1 (n_362), .B2 (n_355));
INV_X1 i_16 (.ZN (n_8), .A (n_9));
AOI21_X1 i_15 (.ZN (n_7), .A (n_360), .B1 (n_354), .B2 (n_8));
AOI21_X1 i_14 (.ZN (n_6), .A (n_360), .B1 (p_0[5]), .B2 (adder[5]));
OAI22_X1 i_13 (.ZN (n_5), .A1 (p_0[6]), .A2 (adder[6]), .B1 (n_350), .B2 (n_7));
XNOR2_X1 i_12 (.ZN (p_1[7]), .A (n_11), .B (n_5));
NOR2_X1 i_11 (.ZN (n_4), .A1 (n_359), .A2 (n_350));
XOR2_X1 i_10 (.Z (p_1[6]), .A (n_7), .B (n_4));
XOR2_X1 i_9 (.Z (p_1[5]), .A (n_9), .B (n_6));
XOR2_X1 i_8 (.Z (p_1[4]), .A (n_362), .B (n_10));
OAI21_X1 i_7 (.ZN (n_3), .A (n_371), .B1 (n_376), .B2 (n_373));
XOR2_X1 i_6 (.Z (p_1[3]), .A (n_364), .B (n_3));
OAI21_X1 i_5 (.ZN (n_2), .A (n_370), .B1 (p_0[2]), .B2 (adder[2]));
XNOR2_X1 i_4 (.ZN (p_1[2]), .A (n_365), .B (n_2));
OAI21_X1 i_3 (.ZN (n_1), .A (n_366), .B1 (p_0[1]), .B2 (adder[1]));
XOR2_X1 i_2 (.Z (p_1[1]), .A (n_367), .B (n_1));
OAI21_X1 i_1 (.ZN (n_0), .A (n_367), .B1 (p_0[0]), .B2 (adder[0]));
INV_X1 i_0 (.ZN (p_1[0]), .A (n_0));

endmodule //datapath__0_16

module datapath (p_0, op1);

output [31:0] p_0;
input [31:0] op1;
wire n_29;
wire n_0;
wire n_28;
wire n_27;
wire n_26;
wire n_1;
wire n_25;
wire n_24;
wire n_2;
wire n_23;
wire n_22;
wire n_21;
wire n_20;
wire n_19;
wire n_18;
wire n_3;
wire n_17;
wire n_16;
wire n_15;
wire n_14;
wire n_13;
wire n_12;
wire n_11;
wire n_10;
wire n_9;
wire n_8;
wire n_4;
wire n_7;
wire n_6;
wire n_5;
wire n_33;
wire n_32;
wire n_31;
wire n_30;


INV_X1 i_64 (.ZN (n_33), .A (op1[25]));
INV_X1 i_63 (.ZN (n_32), .A (op1[21]));
INV_X1 i_62 (.ZN (n_31), .A (op1[14]));
INV_X1 i_61 (.ZN (n_30), .A (op1[11]));
OR3_X1 i_60 (.ZN (n_29), .A1 (op1[2]), .A2 (op1[1]), .A3 (op1[0]));
OR2_X1 i_59 (.ZN (n_28), .A1 (n_29), .A2 (op1[3]));
OR2_X1 i_58 (.ZN (n_27), .A1 (n_28), .A2 (op1[4]));
OR3_X1 i_57 (.ZN (n_26), .A1 (n_27), .A2 (op1[5]), .A3 (op1[6]));
OR2_X1 i_56 (.ZN (n_25), .A1 (n_26), .A2 (op1[7]));
OR3_X1 i_55 (.ZN (n_24), .A1 (n_25), .A2 (op1[8]), .A3 (op1[9]));
NOR2_X1 i_54 (.ZN (n_23), .A1 (n_24), .A2 (op1[10]));
NAND2_X1 i_53 (.ZN (n_22), .A1 (n_23), .A2 (n_30));
NOR2_X1 i_52 (.ZN (n_21), .A1 (n_22), .A2 (op1[12]));
NOR3_X1 i_51 (.ZN (n_20), .A1 (n_22), .A2 (op1[12]), .A3 (op1[13]));
NAND2_X1 i_50 (.ZN (n_19), .A1 (n_20), .A2 (n_31));
OR3_X1 i_49 (.ZN (n_18), .A1 (n_19), .A2 (op1[15]), .A3 (op1[16]));
OR2_X1 i_48 (.ZN (n_17), .A1 (n_18), .A2 (op1[17]));
NOR2_X1 i_47 (.ZN (n_16), .A1 (n_17), .A2 (op1[18]));
NOR3_X1 i_46 (.ZN (n_15), .A1 (n_17), .A2 (op1[18]), .A3 (op1[19]));
NOR4_X1 i_45 (.ZN (n_14), .A1 (n_17), .A2 (op1[18]), .A3 (op1[19]), .A4 (op1[20]));
NAND2_X1 i_44 (.ZN (n_13), .A1 (n_14), .A2 (n_32));
OR2_X1 i_43 (.ZN (n_12), .A1 (n_13), .A2 (op1[22]));
NOR2_X1 i_42 (.ZN (n_11), .A1 (n_12), .A2 (op1[23]));
NOR3_X1 i_41 (.ZN (n_10), .A1 (n_12), .A2 (op1[23]), .A3 (op1[24]));
NAND2_X1 i_40 (.ZN (n_9), .A1 (n_10), .A2 (n_33));
OR3_X1 i_39 (.ZN (n_8), .A1 (n_9), .A2 (op1[26]), .A3 (op1[27]));
NOR2_X1 i_38 (.ZN (n_7), .A1 (n_8), .A2 (op1[28]));
NOR3_X1 i_37 (.ZN (n_6), .A1 (n_8), .A2 (op1[28]), .A3 (op1[29]));
NOR4_X1 i_36 (.ZN (n_5), .A1 (n_8), .A2 (op1[28]), .A3 (op1[29]), .A4 (op1[30]));
XNOR2_X1 i_35 (.ZN (p_0[31]), .A (op1[31]), .B (n_5));
XNOR2_X1 i_34 (.ZN (p_0[30]), .A (op1[30]), .B (n_6));
XNOR2_X1 i_33 (.ZN (p_0[29]), .A (op1[29]), .B (n_7));
XOR2_X1 i_32 (.Z (p_0[28]), .A (op1[28]), .B (n_8));
OAI21_X1 i_31 (.ZN (n_4), .A (op1[27]), .B1 (n_9), .B2 (op1[26]));
AND2_X1 i_30 (.ZN (p_0[27]), .A1 (n_8), .A2 (n_4));
XOR2_X1 i_29 (.Z (p_0[26]), .A (op1[26]), .B (n_9));
XNOR2_X1 i_28 (.ZN (p_0[25]), .A (op1[25]), .B (n_10));
XNOR2_X1 i_27 (.ZN (p_0[24]), .A (op1[24]), .B (n_11));
XOR2_X1 i_26 (.Z (p_0[23]), .A (op1[23]), .B (n_12));
XOR2_X1 i_25 (.Z (p_0[22]), .A (op1[22]), .B (n_13));
XNOR2_X1 i_24 (.ZN (p_0[21]), .A (op1[21]), .B (n_14));
XNOR2_X1 i_23 (.ZN (p_0[20]), .A (op1[20]), .B (n_15));
XNOR2_X1 i_22 (.ZN (p_0[19]), .A (op1[19]), .B (n_16));
XOR2_X1 i_21 (.Z (p_0[18]), .A (op1[18]), .B (n_17));
XOR2_X1 i_20 (.Z (p_0[17]), .A (op1[17]), .B (n_18));
OAI21_X1 i_19 (.ZN (n_3), .A (op1[16]), .B1 (n_19), .B2 (op1[15]));
AND2_X1 i_18 (.ZN (p_0[16]), .A1 (n_18), .A2 (n_3));
XOR2_X1 i_17 (.Z (p_0[15]), .A (op1[15]), .B (n_19));
XNOR2_X1 i_16 (.ZN (p_0[14]), .A (op1[14]), .B (n_20));
XNOR2_X1 i_15 (.ZN (p_0[13]), .A (op1[13]), .B (n_21));
XOR2_X1 i_14 (.Z (p_0[12]), .A (op1[12]), .B (n_22));
XNOR2_X1 i_13 (.ZN (p_0[11]), .A (op1[11]), .B (n_23));
XOR2_X1 i_12 (.Z (p_0[10]), .A (op1[10]), .B (n_24));
OAI21_X1 i_11 (.ZN (n_2), .A (op1[9]), .B1 (n_25), .B2 (op1[8]));
AND2_X1 i_10 (.ZN (p_0[9]), .A1 (n_24), .A2 (n_2));
XOR2_X1 i_9 (.Z (p_0[8]), .A (op1[8]), .B (n_25));
XOR2_X1 i_8 (.Z (p_0[7]), .A (op1[7]), .B (n_26));
OAI21_X1 i_7 (.ZN (n_1), .A (op1[6]), .B1 (n_27), .B2 (op1[5]));
AND2_X1 i_6 (.ZN (p_0[6]), .A1 (n_26), .A2 (n_1));
XOR2_X1 i_5 (.Z (p_0[5]), .A (op1[5]), .B (n_27));
XOR2_X1 i_4 (.Z (p_0[4]), .A (op1[4]), .B (n_28));
XOR2_X1 i_3 (.Z (p_0[3]), .A (op1[3]), .B (n_29));
OAI21_X1 i_2 (.ZN (n_0), .A (op1[2]), .B1 (op1[1]), .B2 (op1[0]));
AND2_X1 i_1 (.ZN (p_0[2]), .A1 (n_29), .A2 (n_0));
XOR2_X1 i_0 (.Z (p_0[1]), .A (op1[1]), .B (op1[0]));

endmodule //datapath

module Radix4_Booth_new (clk, rst, op1, op2, P);

output [63:0] P;
input clk;
input [31:0] op1;
input [31:0] op2;
input rst;
wire n_0_0;
wire n_0_3;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_151;
wire n_0_152;
wire n_0_153;
wire n_0_154;
wire n_0_155;
wire n_0_156;
wire n_0_157;
wire n_0_158;
wire n_0_159;
wire n_0_160;
wire n_0_161;
wire n_0_162;
wire n_0_163;
wire n_0_164;
wire n_0_165;
wire n_0_166;
wire n_0_167;
wire n_0_168;
wire n_0_169;
wire n_0_170;
wire n_0_171;
wire n_0_172;
wire n_0_173;
wire n_0_174;
wire n_0_175;
wire n_0_176;
wire n_0_177;
wire n_0_178;
wire n_0_179;
wire n_0_180;
wire n_0_181;
wire n_0_182;
wire n_0_183;
wire n_0_184;
wire n_0_185;
wire n_0_186;
wire n_0_187;
wire n_0_188;
wire n_0_189;
wire n_0_190;
wire n_0_191;
wire n_0_192;
wire n_0_193;
wire n_0_194;
wire n_0_195;
wire n_0_196;
wire n_0_197;
wire n_0_198;
wire n_0_199;
wire n_0_200;
wire n_0_201;
wire n_0_202;
wire n_0_203;
wire n_0_204;
wire n_0_205;
wire n_0_206;
wire n_0_207;
wire n_0_208;
wire n_0_209;
wire n_0_210;
wire n_0_211;
wire n_0_212;
wire n_0_213;
wire n_0_214;
wire n_0_0_4;
wire n_0_0_0;
wire n_0_0_5;
wire n_0_0_1;
wire n_0_0_6;
wire n_0_0_2;
wire n_0_0_7;
wire n_0_0_3;
wire n_0_279;
wire n_0_280;
wire n_0_281;
wire n_0_282;
wire n_0_283;
wire n_0_284;
wire n_0_285;
wire n_0_286;
wire n_0_287;
wire n_0_288;
wire n_0_289;
wire n_0_290;
wire n_0_291;
wire n_0_292;
wire n_0_293;
wire n_0_294;
wire n_0_295;
wire n_0_296;
wire n_0_1;
wire n_0_2;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_68;
wire n_0_69;
wire n_0_70;
wire n_0_71;
wire n_0_72;
wire n_0_73;
wire n_0_74;
wire n_0_75;
wire n_0_76;
wire n_0_77;
wire n_0_215;
wire n_0_216;
wire n_0_217;
wire n_0_218;
wire n_0_219;
wire n_0_220;
wire n_0_221;
wire n_0_222;
wire n_0_223;
wire n_0_224;
wire n_0_225;
wire n_0_226;
wire n_0_227;
wire n_0_228;
wire n_0_229;
wire n_0_230;
wire n_0_231;
wire n_0_232;
wire n_0_233;
wire n_0_234;
wire n_0_235;
wire n_0_236;
wire n_0_237;
wire n_0_238;
wire n_0_239;
wire n_0_240;
wire n_0_241;
wire n_0_242;
wire n_0_243;
wire n_0_244;
wire n_0_245;
wire n_0_246;
wire n_0_247;
wire n_0_248;
wire n_0_249;
wire n_0_250;
wire n_0_251;
wire n_0_252;
wire n_0_253;
wire n_0_254;
wire n_0_255;
wire n_0_256;
wire n_0_257;
wire n_0_258;
wire n_0_259;
wire n_0_260;
wire n_0_261;
wire n_0_262;
wire n_0_263;
wire n_0_264;
wire n_0_265;
wire n_0_266;
wire n_0_267;
wire n_0_268;
wire n_0_269;
wire n_0_270;
wire n_0_271;
wire n_0_272;
wire n_0_273;
wire n_0_274;
wire n_0_275;
wire n_0_276;
wire n_0_277;
wire n_0_278;
wire n_0_78;
wire n_0_79;
wire n_0_81;
wire n_0_82;
wire n_0_83;
wire n_0_0_8;
wire n_0_84;
wire n_0_85;
wire n_0_0_9;
wire n_0_0_10;
wire n_0_0_11;
wire n_0_0_12;
wire n_0_0_13;
wire n_0_0_14;
wire n_0_0_15;
wire n_0_0_16;
wire n_0_0_17;
wire n_0_0_18;
wire n_0_0_19;
wire n_0_0_20;
wire n_0_80;
wire n_0_86;
wire n_0_90;
wire n_0_91;
wire n_0_92;
wire n_0_0_21;
wire n_0_93;
wire n_0_0_22;
wire n_0_0_23;
wire n_0_94;
wire n_0_0_24;
wire n_0_95;
wire n_0_0_25;
wire n_0_96;
wire n_0_0_26;
wire n_0_0_27;
wire n_0_0_28;
wire n_0_97;
wire n_0_0_29;
wire n_0_98;
wire n_0_0_30;
wire n_0_99;
wire n_0_0_31;
wire n_0_100;
wire n_0_0_32;
wire n_0_101;
wire n_0_0_33;
wire n_0_102;
wire n_0_0_34;
wire n_0_103;
wire n_0_0_35;
wire n_0_0_36;
wire n_0_104;
wire n_0_0_37;
wire n_0_0_38;
wire n_0_105;
wire n_0_0_39;
wire n_0_106;
wire n_0_0_40;
wire n_0_0_41;
wire n_0_107;
wire n_0_0_42;
wire n_0_108;
wire n_0_0_43;
wire n_0_0_44;
wire n_0_0_45;
wire n_0_0_46;
wire n_0_109;
wire n_0_0_47;
wire n_0_110;
wire n_0_0_48;
wire n_0_0_49;
wire n_0_111;
wire n_0_0_50;
wire n_0_0_51;
wire n_0_0_52;
wire n_0_112;
wire n_0_0_53;
wire n_0_0_54;
wire n_0_0_55;
wire n_0_113;
wire n_0_0_56;
wire n_0_0_57;
wire n_0_0_58;
wire n_0_0_59;
wire n_0_0_60;
wire n_0_114;
wire n_0_0_61;
wire n_0_0_62;
wire n_0_0_63;
wire n_0_0_64;
wire n_0_115;
wire n_0_0_65;
wire n_0_0_66;
wire n_0_0_67;
wire n_0_0_68;
wire n_0_0_69;
wire n_0_116;
wire n_0_0_70;
wire n_0_0_71;
wire n_0_0_72;
wire n_0_117;
wire n_0_0_73;
wire n_0_0_74;
wire n_0_0_75;
wire n_0_118;
wire n_0_0_76;
wire n_0_0_77;
wire n_0_0_78;
wire n_0_0_79;
wire n_0_119;
wire n_0_0_80;
wire n_0_0_81;
wire n_0_0_82;
wire n_0_120;
wire n_0_0_83;
wire n_0_0_84;
wire n_0_0_85;
wire n_0_0_86;
wire n_0_0_87;
wire n_0_0_88;
wire n_0_0_89;
wire n_0_0_90;
wire n_0_121;
wire n_0_0_91;
wire n_0_0_92;
wire n_0_0_93;
wire n_0_0_94;
wire n_0_0_95;
wire n_0_0_96;
wire n_0_0_97;
wire n_0_0_98;
wire n_0_122;
wire n_0_0_99;
wire n_0_0_100;
wire n_0_0_101;
wire n_0_0_102;
wire n_0_0_103;
wire n_0_0_104;
wire n_0_0_105;
wire n_0_123;
wire n_0_0_106;
wire n_0_0_107;
wire n_0_0_108;
wire n_0_0_109;
wire n_0_0_110;
wire n_0_0_111;
wire n_0_0_112;
wire n_0_0_113;
wire n_0_0_114;
wire n_0_124;
wire n_0_0_115;
wire n_0_0_116;
wire n_0_0_117;
wire n_0_0_118;
wire n_0_0_119;
wire n_0_0_120;
wire n_0_0_121;
wire n_0_0_122;
wire n_0_125;
wire n_0_0_123;
wire n_0_0_124;
wire n_0_0_125;
wire n_0_0_126;
wire n_0_0_127;
wire n_0_0_128;
wire n_0_0_129;
wire n_0_0_130;
wire n_0_0_131;
wire n_0_126;
wire n_0_0_132;
wire n_0_0_133;
wire n_0_0_134;
wire n_0_0_135;
wire n_0_0_136;
wire n_0_0_137;
wire n_0_0_138;
wire n_0_127;
wire n_0_0_139;
wire n_0_0_140;
wire n_0_0_141;
wire n_0_0_142;
wire n_0_0_143;
wire n_0_0_144;
wire n_0_0_145;
wire n_0_128;
wire n_0_0_146;
wire n_0_0_147;
wire n_0_0_148;
wire n_0_0_149;
wire n_0_0_150;
wire n_0_0_151;
wire n_0_0_152;
wire n_0_0_153;
wire n_0_129;
wire n_0_0_154;
wire n_0_0_155;
wire n_0_0_156;
wire n_0_0_157;
wire n_0_0_158;
wire n_0_0_159;
wire n_0_0_160;
wire n_0_130;
wire n_0_0_161;
wire n_0_0_162;
wire n_0_0_163;
wire n_0_0_164;
wire n_0_0_165;
wire n_0_0_166;
wire n_0_131;
wire n_0_0_167;
wire n_0_0_168;
wire n_0_0_169;
wire n_0_0_170;
wire n_0_0_171;
wire n_0_0_172;
wire n_0_0_173;
wire n_0_132;
wire n_0_0_174;
wire n_0_0_175;
wire n_0_0_176;
wire n_0_0_177;
wire n_0_0_178;
wire n_0_0_179;
wire n_0_0_180;
wire n_0_133;
wire n_0_0_181;
wire n_0_0_182;
wire n_0_0_183;
wire n_0_0_184;
wire n_0_0_185;
wire n_0_0_186;
wire n_0_0_187;
wire n_0_134;
wire n_0_0_188;
wire n_0_0_189;
wire n_0_0_190;
wire n_0_0_191;
wire n_0_0_192;
wire n_0_0_193;
wire n_0_0_194;
wire n_0_135;
wire n_0_0_195;
wire n_0_0_196;
wire n_0_0_197;
wire n_0_0_198;
wire n_0_0_199;
wire n_0_0_200;
wire n_0_136;
wire n_0_0_201;
wire n_0_0_202;
wire n_0_0_203;
wire n_0_0_204;
wire n_0_0_205;
wire n_0_0_206;
wire n_0_137;
wire n_0_0_207;
wire n_0_0_208;
wire n_0_0_209;
wire n_0_0_210;
wire n_0_0_211;
wire n_0_0_212;
wire n_0_0_213;
wire n_0_138;
wire n_0_0_214;
wire n_0_0_215;
wire n_0_0_216;
wire n_0_0_217;
wire n_0_0_218;
wire n_0_0_219;
wire n_0_0_220;
wire n_0_139;
wire n_0_0_221;
wire n_0_0_222;
wire n_0_0_223;
wire n_0_0_224;
wire n_0_0_225;
wire n_0_0_226;
wire n_0_0_227;
wire n_0_140;
wire n_0_0_228;
wire n_0_0_229;
wire n_0_0_230;
wire n_0_0_231;
wire n_0_0_232;
wire n_0_0_233;
wire n_0_0_234;
wire n_0_141;
wire n_0_0_235;
wire n_0_0_236;
wire n_0_0_237;
wire n_0_0_238;
wire n_0_0_239;
wire n_0_0_240;
wire n_0_142;
wire n_0_0_241;
wire n_0_0_242;
wire n_0_0_243;
wire n_0_0_244;
wire n_0_0_245;
wire n_0_0_246;
wire n_0_0_247;
wire n_0_0_248;
wire n_0_143;
wire n_0_0_249;
wire n_0_0_250;
wire n_0_0_251;
wire n_0_0_252;
wire n_0_0_253;
wire n_0_0_254;
wire n_0_144;
wire n_0_0_255;
wire n_0_0_256;
wire n_0_0_257;
wire n_0_0_258;
wire n_0_0_259;
wire n_0_145;
wire n_0_0_260;
wire n_0_0_261;
wire n_0_0_262;
wire n_0_0_263;
wire n_0_0_264;
wire n_0_0_265;
wire n_0_146;
wire n_0_0_266;
wire n_0_0_267;
wire n_0_0_268;
wire n_0_0_269;
wire n_0_0_270;
wire n_0_0_271;
wire n_0_147;
wire n_0_0_272;
wire n_0_0_273;
wire n_0_0_274;
wire n_0_0_275;
wire n_0_0_276;
wire n_0_0_277;
wire n_0_148;
wire n_0_0_278;
wire n_0_0_279;
wire n_0_0_280;
wire n_0_0_281;
wire n_0_0_282;
wire n_0_0_283;
wire n_0_149;
wire n_0_0_284;
wire n_0_0_285;
wire n_0_0_286;
wire n_0_0_287;
wire n_0_0_288;
wire n_0_0_289;
wire n_0_150;
wire n_0_0_290;
wire n_0_0_291;
wire n_0_0_292;
wire n_0_0_293;
wire n_0_0_294;
wire n_0_0_295;
wire n_0_0_296;
wire n_0_0_297;
wire n_0_0_298;
wire n_0_0_299;
wire n_0_89;
wire n_0_0_300;
wire n_0_0_301;
wire n_0_0_302;
wire n_0_0_303;
wire n_0_0_304;
wire n_0_0_305;
wire n_0_0_306;
wire n_0_0_307;
wire n_0_0_308;
wire n_0_0_309;
wire n_0_0_310;
wire n_0_0_311;
wire n_0_0_312;
wire n_0_0_313;
wire n_0_0_314;
wire n_0_0_315;
wire n_0_0_316;
wire n_0_0_317;
wire n_0_0_318;
wire n_0_0_319;
wire n_0_0_320;
wire n_0_0_321;
wire n_0_0_322;
wire n_0_0_323;
wire n_0_0_324;
wire n_0_0_325;
wire n_0_0_326;
wire n_0_0_327;
wire n_0_0_328;
wire n_0_0_329;
wire n_0_0_330;
wire n_0_0_331;
wire n_0_0_332;
wire n_0_0_333;
wire n_0_0_334;
wire n_0_0_335;
wire n_0_0_336;
wire n_0_0_337;
wire n_0_0_338;
wire n_0_0_339;
wire n_0_0_340;
wire n_0_0_341;
wire n_0_0_342;
wire n_0_0_343;
wire n_0_0_344;
wire n_0_0_345;
wire n_0_0_346;
wire n_0_0_347;
wire n_0_0_348;
wire n_0_0_349;
wire n_0_0_350;
wire n_0_0_351;
wire n_0_0_352;
wire n_0_0_353;
wire n_0_0_354;
wire n_0_0_355;
wire n_0_0_356;
wire n_0_0_357;
wire n_0_0_358;
wire n_0_0_359;
wire \adder[63] ;
wire \adder[62] ;
wire \adder[61] ;
wire \adder[60] ;
wire \adder[59] ;
wire \adder[58] ;
wire \adder[57] ;
wire \adder[56] ;
wire \adder[55] ;
wire \adder[54] ;
wire \adder[53] ;
wire \adder[52] ;
wire \adder[51] ;
wire \adder[50] ;
wire \adder[49] ;
wire \adder[48] ;
wire \adder[47] ;
wire \adder[46] ;
wire \adder[45] ;
wire \adder[44] ;
wire \adder[43] ;
wire \adder[42] ;
wire \adder[41] ;
wire \adder[40] ;
wire \adder[39] ;
wire \adder[38] ;
wire \adder[37] ;
wire \adder[36] ;
wire \adder[35] ;
wire \adder[34] ;
wire \adder[33] ;
wire \adder[32] ;
wire \adder[31] ;
wire \adder[30] ;
wire \adder[29] ;
wire \adder[28] ;
wire \adder[27] ;
wire \adder[26] ;
wire \adder[25] ;
wire \adder[24] ;
wire \adder[23] ;
wire \adder[22] ;
wire \adder[21] ;
wire \adder[20] ;
wire \adder[19] ;
wire \adder[18] ;
wire \adder[17] ;
wire \adder[16] ;
wire \adder[15] ;
wire \adder[14] ;
wire \adder[13] ;
wire \adder[12] ;
wire \adder[11] ;
wire \adder[10] ;
wire \adder[9] ;
wire \adder[8] ;
wire \adder[7] ;
wire \adder[6] ;
wire \adder[5] ;
wire \adder[4] ;
wire \adder[3] ;
wire \adder[2] ;
wire \adder[1] ;
wire \adder[0] ;
wire \n[5] ;
wire \n[4] ;
wire \n[3] ;
wire \n[2] ;
wire \n[1] ;
wire \n[0] ;
wire n_0_87;
wire \OP1_complement[31] ;
wire \OP1_complement[30] ;
wire \OP1_complement[29] ;
wire \OP1_complement[28] ;
wire \OP1_complement[27] ;
wire \OP1_complement[26] ;
wire \OP1_complement[25] ;
wire \OP1_complement[24] ;
wire \OP1_complement[23] ;
wire \OP1_complement[22] ;
wire \OP1_complement[21] ;
wire \OP1_complement[20] ;
wire \OP1_complement[19] ;
wire \OP1_complement[18] ;
wire \OP1_complement[17] ;
wire \OP1_complement[16] ;
wire \OP1_complement[15] ;
wire \OP1_complement[14] ;
wire \OP1_complement[13] ;
wire \OP1_complement[12] ;
wire \OP1_complement[11] ;
wire \OP1_complement[10] ;
wire \OP1_complement[9] ;
wire \OP1_complement[8] ;
wire \OP1_complement[7] ;
wire \OP1_complement[6] ;
wire \OP1_complement[5] ;
wire \OP1_complement[4] ;
wire \OP1_complement[3] ;
wire \OP1_complement[2] ;
wire \OP1_complement[1] ;
wire \OP1_complement[0] ;
wire q;
wire n_0_88;
wire uc_0;
wire uc_1;
wire uc_2;
wire sps__n1;
wire sps__n4;
wire sps__n7;
wire sps__n10;
wire sps__n11;
wire sps__n16;
wire spc__n19;
wire spc__n22;
wire spt__n25;


CLKGATETST_X1 clk_gate_adder_reg (.GCK (n_0_88), .CK (clk), .E (n_0_84), .SE (1'b0 ));
DFF_X1 q_reg (.Q (q), .CK (n_0_88), .D (n_0_85));
DFF_X1 \OP1_complement_reg[0]  (.Q (\OP1_complement[0] ), .CK (n_0_87), .D (op1[0]));
DFF_X1 \OP1_complement_reg[1]  (.Q (\OP1_complement[1] ), .CK (n_0_87), .D (n_0_3));
DFF_X1 \OP1_complement_reg[2]  (.Q (\OP1_complement[2] ), .CK (n_0_87), .D (n_0_4));
DFF_X1 \OP1_complement_reg[3]  (.Q (\OP1_complement[3] ), .CK (n_0_87), .D (n_0_5));
DFF_X1 \OP1_complement_reg[4]  (.Q (\OP1_complement[4] ), .CK (n_0_87), .D (n_0_6));
DFF_X1 \OP1_complement_reg[5]  (.Q (\OP1_complement[5] ), .CK (n_0_87), .D (n_0_7));
DFF_X1 \OP1_complement_reg[6]  (.Q (\OP1_complement[6] ), .CK (n_0_87), .D (n_0_8));
DFF_X1 \OP1_complement_reg[7]  (.Q (\OP1_complement[7] ), .CK (n_0_87), .D (n_0_9));
DFF_X1 \OP1_complement_reg[8]  (.Q (\OP1_complement[8] ), .CK (n_0_87), .D (n_0_10));
DFF_X1 \OP1_complement_reg[9]  (.Q (\OP1_complement[9] ), .CK (n_0_87), .D (n_0_11));
DFF_X1 \OP1_complement_reg[10]  (.Q (\OP1_complement[10] ), .CK (n_0_87), .D (n_0_12));
DFF_X1 \OP1_complement_reg[11]  (.Q (\OP1_complement[11] ), .CK (n_0_87), .D (n_0_13));
DFF_X1 \OP1_complement_reg[12]  (.Q (\OP1_complement[12] ), .CK (n_0_87), .D (n_0_14));
DFF_X1 \OP1_complement_reg[13]  (.Q (\OP1_complement[13] ), .CK (n_0_87), .D (n_0_15));
DFF_X1 \OP1_complement_reg[14]  (.Q (\OP1_complement[14] ), .CK (n_0_87), .D (n_0_16));
DFF_X1 \OP1_complement_reg[15]  (.Q (\OP1_complement[15] ), .CK (n_0_87), .D (n_0_17));
DFF_X1 \OP1_complement_reg[16]  (.Q (\OP1_complement[16] ), .CK (n_0_87), .D (n_0_18));
DFF_X1 \OP1_complement_reg[17]  (.Q (\OP1_complement[17] ), .CK (n_0_87), .D (n_0_19));
DFF_X1 \OP1_complement_reg[18]  (.Q (\OP1_complement[18] ), .CK (n_0_87), .D (n_0_20));
DFF_X1 \OP1_complement_reg[19]  (.Q (\OP1_complement[19] ), .CK (n_0_87), .D (n_0_21));
DFF_X1 \OP1_complement_reg[20]  (.Q (\OP1_complement[20] ), .CK (n_0_87), .D (n_0_22));
DFF_X1 \OP1_complement_reg[21]  (.Q (\OP1_complement[21] ), .CK (n_0_87), .D (n_0_23));
DFF_X1 \OP1_complement_reg[22]  (.Q (\OP1_complement[22] ), .CK (n_0_87), .D (n_0_24));
DFF_X1 \OP1_complement_reg[23]  (.Q (\OP1_complement[23] ), .CK (n_0_87), .D (n_0_25));
DFF_X1 \OP1_complement_reg[24]  (.Q (\OP1_complement[24] ), .CK (n_0_87), .D (n_0_26));
DFF_X1 \OP1_complement_reg[25]  (.Q (\OP1_complement[25] ), .CK (n_0_87), .D (n_0_27));
DFF_X1 \OP1_complement_reg[26]  (.Q (\OP1_complement[26] ), .CK (n_0_87), .D (n_0_28));
DFF_X1 \OP1_complement_reg[27]  (.Q (\OP1_complement[27] ), .CK (n_0_87), .D (n_0_29));
DFF_X1 \OP1_complement_reg[28]  (.Q (\OP1_complement[28] ), .CK (n_0_87), .D (n_0_30));
DFF_X1 \OP1_complement_reg[29]  (.Q (\OP1_complement[29] ), .CK (n_0_87), .D (n_0_31));
DFF_X1 \OP1_complement_reg[30]  (.Q (\OP1_complement[30] ), .CK (n_0_87), .D (n_0_32));
DFF_X1 \OP1_complement_reg[31]  (.Q (\OP1_complement[31] ), .CK (n_0_87), .D (n_0_33));
CLKGATETST_X1 clk_gate_OP1_complement_reg (.GCK (n_0_87), .CK (clk), .E (rst), .SE (1'b0 ));
DFF_X1 \n_reg[0]  (.Q (\n[0] ), .CK (n_0_88), .D (n_0_78));
DFF_X1 \n_reg[1]  (.Q (\n[1] ), .CK (n_0_88), .D (n_0_79));
DFF_X1 \n_reg[2]  (.Q (spt__n25), .CK (n_0_88), .D (n_0_80));
DFF_X1 \n_reg[3]  (.Q (\n[3] ), .CK (n_0_88), .D (n_0_81));
DFF_X1 \n_reg[4]  (.Q (\n[4] ), .CK (n_0_88), .D (n_0_82));
DFF_X1 \n_reg[5]  (.Q (\n[5] ), .CK (n_0_88), .D (n_0_83));
DFF_X1 \adder_reg[0]  (.Q (\adder[0] ), .CK (n_0_88), .D (n_0_215));
DFF_X1 \adder_reg[1]  (.Q (\adder[1] ), .CK (n_0_88), .D (n_0_216));
DFF_X1 \adder_reg[2]  (.Q (\adder[2] ), .CK (n_0_88), .D (n_0_217));
DFF_X1 \adder_reg[3]  (.Q (\adder[3] ), .CK (n_0_88), .D (n_0_218));
DFF_X1 \adder_reg[4]  (.Q (\adder[4] ), .CK (n_0_88), .D (n_0_219));
DFF_X1 \adder_reg[5]  (.Q (\adder[5] ), .CK (n_0_88), .D (n_0_220));
DFF_X1 \adder_reg[6]  (.Q (\adder[6] ), .CK (n_0_88), .D (n_0_221));
DFF_X1 \adder_reg[7]  (.Q (\adder[7] ), .CK (n_0_88), .D (n_0_222));
DFF_X1 \adder_reg[8]  (.Q (\adder[8] ), .CK (n_0_88), .D (n_0_223));
DFF_X1 \adder_reg[9]  (.Q (\adder[9] ), .CK (n_0_88), .D (n_0_224));
DFF_X1 \adder_reg[10]  (.Q (\adder[10] ), .CK (n_0_88), .D (n_0_225));
DFF_X1 \adder_reg[11]  (.Q (\adder[11] ), .CK (n_0_88), .D (n_0_226));
DFF_X1 \adder_reg[12]  (.Q (\adder[12] ), .CK (n_0_88), .D (n_0_227));
DFF_X1 \adder_reg[13]  (.Q (\adder[13] ), .CK (n_0_88), .D (n_0_228));
DFF_X1 \adder_reg[14]  (.Q (\adder[14] ), .CK (n_0_88), .D (n_0_229));
DFF_X1 \adder_reg[15]  (.Q (\adder[15] ), .CK (n_0_88), .D (n_0_230));
DFF_X1 \adder_reg[16]  (.Q (\adder[16] ), .CK (n_0_88), .D (n_0_231));
DFF_X1 \adder_reg[17]  (.Q (\adder[17] ), .CK (n_0_88), .D (n_0_232));
DFF_X1 \adder_reg[18]  (.Q (\adder[18] ), .CK (n_0_88), .D (n_0_233));
DFF_X1 \adder_reg[19]  (.Q (\adder[19] ), .CK (n_0_88), .D (n_0_234));
DFF_X1 \adder_reg[20]  (.Q (\adder[20] ), .CK (n_0_88), .D (n_0_235));
DFF_X1 \adder_reg[21]  (.Q (\adder[21] ), .CK (n_0_88), .D (n_0_236));
DFF_X1 \adder_reg[22]  (.Q (\adder[22] ), .CK (n_0_88), .D (n_0_237));
DFF_X1 \adder_reg[23]  (.Q (\adder[23] ), .CK (n_0_88), .D (n_0_238));
DFF_X1 \adder_reg[24]  (.Q (\adder[24] ), .CK (n_0_88), .D (n_0_239));
DFF_X1 \adder_reg[25]  (.Q (\adder[25] ), .CK (n_0_88), .D (n_0_240));
DFF_X1 \adder_reg[26]  (.Q (\adder[26] ), .CK (n_0_88), .D (n_0_241));
DFF_X1 \adder_reg[27]  (.Q (\adder[27] ), .CK (n_0_88), .D (n_0_242));
DFF_X1 \adder_reg[28]  (.Q (\adder[28] ), .CK (n_0_88), .D (n_0_243));
DFF_X1 \adder_reg[29]  (.Q (\adder[29] ), .CK (n_0_88), .D (n_0_244));
DFF_X1 \adder_reg[30]  (.Q (\adder[30] ), .CK (n_0_88), .D (n_0_245));
DFF_X1 \adder_reg[31]  (.Q (\adder[31] ), .CK (n_0_88), .D (n_0_246));
DFF_X1 \adder_reg[32]  (.Q (\adder[32] ), .CK (n_0_88), .D (n_0_247));
DFF_X1 \adder_reg[33]  (.Q (\adder[33] ), .CK (n_0_88), .D (n_0_248));
DFF_X1 \adder_reg[34]  (.Q (\adder[34] ), .CK (n_0_88), .D (n_0_249));
DFF_X1 \adder_reg[35]  (.Q (\adder[35] ), .CK (n_0_88), .D (n_0_250));
DFF_X1 \adder_reg[36]  (.Q (\adder[36] ), .CK (n_0_88), .D (n_0_251));
DFF_X1 \adder_reg[37]  (.Q (\adder[37] ), .CK (n_0_88), .D (n_0_252));
DFF_X1 \adder_reg[38]  (.Q (\adder[38] ), .CK (n_0_88), .D (n_0_253));
DFF_X1 \adder_reg[39]  (.Q (\adder[39] ), .CK (n_0_88), .D (n_0_254));
DFF_X1 \adder_reg[40]  (.Q (\adder[40] ), .CK (n_0_88), .D (n_0_255));
DFF_X1 \adder_reg[41]  (.Q (\adder[41] ), .CK (n_0_88), .D (n_0_256));
DFF_X1 \adder_reg[42]  (.Q (\adder[42] ), .CK (n_0_88), .D (n_0_257));
DFF_X1 \adder_reg[43]  (.Q (\adder[43] ), .CK (n_0_88), .D (n_0_258));
DFF_X1 \adder_reg[44]  (.Q (\adder[44] ), .CK (n_0_88), .D (n_0_259));
DFF_X1 \adder_reg[45]  (.Q (\adder[45] ), .CK (n_0_88), .D (n_0_260));
DFF_X1 \adder_reg[46]  (.Q (\adder[46] ), .CK (n_0_88), .D (n_0_261));
DFF_X1 \adder_reg[47]  (.Q (\adder[47] ), .CK (n_0_88), .D (n_0_262));
DFF_X1 \adder_reg[48]  (.Q (\adder[48] ), .CK (n_0_88), .D (n_0_263));
DFF_X1 \adder_reg[49]  (.Q (\adder[49] ), .CK (n_0_88), .D (n_0_264));
DFF_X1 \adder_reg[50]  (.Q (\adder[50] ), .CK (n_0_88), .D (n_0_265));
DFF_X1 \adder_reg[51]  (.Q (\adder[51] ), .CK (n_0_88), .D (n_0_266));
DFF_X1 \adder_reg[52]  (.Q (\adder[52] ), .CK (n_0_88), .D (n_0_267));
DFF_X1 \adder_reg[53]  (.Q (\adder[53] ), .CK (n_0_88), .D (n_0_268));
DFF_X1 \adder_reg[54]  (.Q (\adder[54] ), .CK (n_0_88), .D (n_0_269));
DFF_X1 \adder_reg[55]  (.Q (\adder[55] ), .CK (n_0_88), .D (n_0_270));
DFF_X1 \adder_reg[56]  (.Q (\adder[56] ), .CK (n_0_88), .D (n_0_271));
DFF_X1 \adder_reg[57]  (.Q (\adder[57] ), .CK (n_0_88), .D (n_0_272));
DFF_X1 \adder_reg[58]  (.Q (\adder[58] ), .CK (n_0_88), .D (n_0_273));
DFF_X1 \adder_reg[59]  (.Q (\adder[59] ), .CK (n_0_88), .D (n_0_274));
DFF_X1 \adder_reg[60]  (.Q (\adder[60] ), .CK (n_0_88), .D (n_0_275));
DFF_X1 \adder_reg[61]  (.Q (\adder[61] ), .CK (n_0_88), .D (n_0_276));
DFF_X1 \adder_reg[62]  (.Q (\adder[62] ), .CK (n_0_88), .D (n_0_277));
DFF_X1 \adder_reg[63]  (.Q (\adder[63] ), .CK (n_0_88), .D (n_0_278));
INV_X1 i_0_0_554 (.ZN (n_0_0_359), .A (\n[3] ));
INV_X1 i_0_0_553 (.ZN (n_0_0_358), .A (\n[2] ));
INV_X1 i_0_0_552 (.ZN (n_0_0_357), .A (sps__n7));
INV_X4 i_0_0_551 (.ZN (n_0_0_356), .A (sps__n11));
INV_X1 i_0_0_550 (.ZN (n_0_0_355), .A (q));
INV_X4 i_0_0_549 (.ZN (n_0_0_354), .A (rst));
INV_X1 i_0_0_548 (.ZN (n_0_0_353), .A (n_0_0_4));
INV_X1 i_0_0_547 (.ZN (n_0_0_352), .A (n_0_0_5));
INV_X1 i_0_0_546 (.ZN (n_0_0_351), .A (n_0_0_6));
NAND2_X1 i_0_0_545 (.ZN (n_0_0_350), .A1 (n_0_0_359), .A2 (\n[2] ));
INV_X1 i_0_0_544 (.ZN (n_0_0_349), .A (n_0_0_350));
NOR3_X1 i_0_0_543 (.ZN (n_0_0_348), .A1 (sps__n7), .A2 (n_0_0_356), .A3 (n_0_0_350));
AOI22_X1 i_0_0_542 (.ZN (n_0_0_347), .A1 (sps__n1), .A2 (op2[8]), .B1 (sps__n7), .B2 (op2[12]));
AOI22_X1 i_0_0_541 (.ZN (n_0_0_346), .A1 (n_0_0_356), .A2 (op2[28]), .B1 (sps__n11), .B2 (op2[30]));
NAND2_X1 i_0_0_540 (.ZN (n_0_0_345), .A1 (\n[3] ), .A2 (\n[2] ));
INV_X1 i_0_0_539 (.ZN (n_0_0_344), .A (n_0_0_345));
NAND2_X2 i_0_0_538 (.ZN (n_0_0_343), .A1 (\n[3] ), .A2 (n_0_0_358));
INV_X1 i_0_0_537 (.ZN (n_0_0_342), .A (n_0_0_343));
AOI22_X1 i_0_0_536 (.ZN (n_0_0_341), .A1 (op2[26]), .A2 (n_0_0_344), .B1 (op2[18]), .B2 (n_0_0_342));
NAND2_X1 i_0_0_535 (.ZN (n_0_0_340), .A1 (n_0_0_359), .A2 (n_0_0_358));
INV_X1 i_0_0_534 (.ZN (n_0_0_339), .A (n_0_0_340));
NOR3_X1 i_0_0_533 (.ZN (n_0_0_338), .A1 (sps__n7), .A2 (n_0_0_356), .A3 (n_0_0_340));
AOI22_X1 i_0_0_532 (.ZN (n_0_0_337), .A1 (sps__n1), .A2 (op2[0]), .B1 (sps__n7), .B2 (op2[4]));
AOI222_X1 i_0_0_531 (.ZN (n_0_0_336), .A1 (op2[6]), .A2 (n_0_0_339), .B1 (op2[22])
    , .B2 (n_0_0_342), .C1 (op2[14]), .C2 (n_0_0_349));
OR3_X1 i_0_0_530 (.ZN (n_0_0_335), .A1 (sps__n1), .A2 (n_0_0_356), .A3 (n_0_0_336));
AOI21_X1 i_0_0_529 (.ZN (n_0_0_334), .A (sps__n1), .B1 (op2[20]), .B2 (n_0_0_342));
AOI221_X1 i_0_0_528 (.ZN (n_0_0_333), .A (sps__n7), .B1 (op2[24]), .B2 (n_0_0_344)
    , .C1 (op2[16]), .C2 (n_0_0_342));
OR3_X1 i_0_0_527 (.ZN (n_0_0_332), .A1 (sps__n11), .A2 (n_0_0_334), .A3 (n_0_0_333));
OAI33_X1 i_0_0_526 (.ZN (n_0_0_331), .A1 (sps__n11), .A2 (n_0_0_350), .A3 (n_0_0_347)
    , .B1 (sps__n11), .B2 (n_0_0_340), .B3 (n_0_0_337));
AOI221_X1 i_0_0_525 (.ZN (n_0_0_330), .A (n_0_0_331), .B1 (op2[10]), .B2 (n_0_0_348)
    , .C1 (op2[2]), .C2 (n_0_0_338));
OAI33_X1 i_0_0_524 (.ZN (n_0_0_329), .A1 (n_0_0_346), .A2 (n_0_0_345), .A3 (sps__n1)
    , .B1 (sps__n7), .B2 (n_0_0_356), .B3 (n_0_0_341));
INV_X1 i_0_0_523 (.ZN (n_0_0_328), .A (n_0_0_329));
NAND4_X1 i_0_0_522 (.ZN (n_0_0_327), .A1 (n_0_0_332), .A2 (n_0_0_330), .A3 (n_0_0_335), .A4 (n_0_0_328));
INV_X1 i_0_0_521 (.ZN (n_0_0_326), .A (n_0_0_327));
AOI22_X1 i_0_0_520 (.ZN (n_0_0_325), .A1 (q), .A2 (n_0_0_327), .B1 (n_0_0_355), .B2 (n_0_0_326));
AOI221_X1 i_0_0_519 (.ZN (n_0_0_324), .A (sps__n7), .B1 (n_0_0_356), .B2 (op2[17])
    , .C1 (sps__n11), .C2 (op2[19]));
AOI221_X1 i_0_0_518 (.ZN (n_0_0_323), .A (sps__n1), .B1 (sps__n11), .B2 (op2[23])
    , .C1 (n_0_0_356), .C2 (op2[21]));
AOI221_X1 i_0_0_517 (.ZN (n_0_0_322), .A (sps__n1), .B1 (sps__n11), .B2 (op2[31])
    , .C1 (n_0_0_356), .C2 (op2[29]));
AOI221_X1 i_0_0_516 (.ZN (n_0_0_321), .A (sps__n7), .B1 (n_0_0_356), .B2 (op2[25])
    , .C1 (sps__n11), .C2 (op2[27]));
OAI33_X1 i_0_0_515 (.ZN (n_0_0_320), .A1 (n_0_0_324), .A2 (n_0_0_323), .A3 (n_0_0_343)
    , .B1 (n_0_0_322), .B2 (n_0_0_321), .B3 (n_0_0_345));
INV_X1 i_0_0_514 (.ZN (n_0_0_319), .A (n_0_0_320));
AOI22_X1 i_0_0_513 (.ZN (n_0_0_318), .A1 (op2[15]), .A2 (n_0_0_349), .B1 (op2[7]), .B2 (n_0_0_339));
OR3_X1 i_0_0_512 (.ZN (n_0_0_317), .A1 (sps__n1), .A2 (n_0_0_356), .A3 (n_0_0_318));
NOR2_X1 i_0_0_511 (.ZN (n_0_0_316), .A1 (\n[3] ), .A2 (sps__n7));
NAND2_X1 i_0_0_510 (.ZN (n_0_0_315), .A1 (n_0_0_358), .A2 (n_0_0_316));
INV_X1 i_0_0_509 (.ZN (n_0_0_314), .A (n_0_0_315));
AOI22_X1 i_0_0_508 (.ZN (n_0_0_313), .A1 (sps__n1), .A2 (op2[9]), .B1 (sps__n7), .B2 (op2[13]));
NOR3_X1 i_0_0_507 (.ZN (n_0_0_312), .A1 (sps__n11), .A2 (n_0_0_350), .A3 (n_0_0_313));
AOI21_X1 i_0_0_506 (.ZN (n_0_0_311), .A (n_0_0_312), .B1 (op2[3]), .B2 (n_0_0_338));
AOI22_X1 i_0_0_505 (.ZN (n_0_0_310), .A1 (sps__n1), .A2 (op2[1]), .B1 (sps__n7), .B2 (op2[5]));
NOR3_X1 i_0_0_504 (.ZN (n_0_0_309), .A1 (sps__n11), .A2 (n_0_0_340), .A3 (n_0_0_310));
AOI21_X1 i_0_0_503 (.ZN (n_0_0_308), .A (n_0_0_309), .B1 (op2[11]), .B2 (n_0_0_348));
NAND4_X1 i_0_0_502 (.ZN (n_0_0_307), .A1 (n_0_0_311), .A2 (n_0_0_308), .A3 (n_0_0_317), .A4 (n_0_0_319));
INV_X1 i_0_0_501 (.ZN (n_0_0_306), .A (n_0_0_307));
AND2_X1 i_0_0_500 (.ZN (n_0_0_305), .A1 (n_0_0_325), .A2 (n_0_0_306));
AND2_X1 i_0_0_499 (.ZN (n_0_0_304), .A1 (n_0_0_325), .A2 (n_0_0_307));
NOR3_X2 i_0_0_498 (.ZN (n_0_0_303), .A1 (n_0_0_355), .A2 (n_0_0_326), .A3 (n_0_0_307));
NOR3_X1 i_0_0_497 (.ZN (n_0_0_302), .A1 (q), .A2 (n_0_0_327), .A3 (n_0_0_306));
AOI22_X1 i_0_0_496 (.ZN (n_0_0_301), .A1 (op1[31]), .A2 (spc__n22), .B1 (\OP1_complement[30] ), .B2 (sps__n16));
AOI22_X1 i_0_0_495 (.ZN (n_0_0_300), .A1 (\OP1_complement[31] ), .A2 (spc__n19), .B1 (op1[30]), .B2 (sps__n4));
NAND2_X1 i_0_0_494 (.ZN (n_0_89), .A1 (n_0_0_301), .A2 (n_0_0_300));
INV_X1 i_0_0_493 (.ZN (n_0_0_299), .A (n_0_89));
NOR2_X1 i_0_0_492 (.ZN (n_0_0_298), .A1 (sps__n11), .A2 (n_0_89));
NOR2_X1 i_0_0_491 (.ZN (n_0_0_297), .A1 (sps__n7), .A2 (n_0_0_299));
NOR2_X1 i_0_0_490 (.ZN (n_0_0_296), .A1 (n_0_0_344), .A2 (n_0_89));
AOI22_X1 i_0_0_489 (.ZN (n_0_0_295), .A1 (op1[30]), .A2 (spc__n22), .B1 (op1[29]), .B2 (sps__n4));
AOI22_X1 i_0_0_488 (.ZN (n_0_0_294), .A1 (\OP1_complement[30] ), .A2 (spc__n19), .B1 (\OP1_complement[29] ), .B2 (sps__n16));
NAND2_X1 i_0_0_487 (.ZN (n_0_0_293), .A1 (n_0_0_295), .A2 (n_0_0_294));
INV_X1 i_0_0_486 (.ZN (n_0_0_292), .A (n_0_0_293));
AOI21_X1 i_0_0_485 (.ZN (n_0_0_291), .A (n_0_0_296), .B1 (n_0_0_344), .B2 (n_0_0_292));
AOI21_X1 i_0_0_484 (.ZN (n_0_0_290), .A (n_0_0_297), .B1 (sps__n7), .B2 (n_0_0_291));
AOI21_X1 i_0_0_483 (.ZN (n_0_150), .A (n_0_0_298), .B1 (sps__n11), .B2 (n_0_0_290));
AOI22_X1 i_0_0_482 (.ZN (n_0_0_289), .A1 (\OP1_complement[29] ), .A2 (spc__n19), .B1 (op1[28]), .B2 (sps__n4));
AOI22_X1 i_0_0_481 (.ZN (n_0_0_288), .A1 (op1[29]), .A2 (spc__n22), .B1 (\OP1_complement[28] ), .B2 (sps__n16));
NAND2_X1 i_0_0_480 (.ZN (n_0_0_287), .A1 (n_0_0_289), .A2 (n_0_0_288));
INV_X1 i_0_0_479 (.ZN (n_0_0_286), .A (n_0_0_287));
AOI21_X1 i_0_0_478 (.ZN (n_0_0_285), .A (n_0_0_296), .B1 (n_0_0_344), .B2 (n_0_0_286));
AOI21_X1 i_0_0_477 (.ZN (n_0_0_284), .A (n_0_0_297), .B1 (sps__n7), .B2 (n_0_0_285));
AOI21_X1 i_0_0_476 (.ZN (n_0_149), .A (n_0_0_298), .B1 (sps__n11), .B2 (n_0_0_284));
AOI22_X1 i_0_0_475 (.ZN (n_0_0_283), .A1 (op1[28]), .A2 (spc__n22), .B1 (\OP1_complement[27] ), .B2 (sps__n16));
AOI22_X1 i_0_0_474 (.ZN (n_0_0_282), .A1 (\OP1_complement[28] ), .A2 (spc__n19), .B1 (op1[27]), .B2 (sps__n4));
NAND2_X1 i_0_0_473 (.ZN (n_0_0_281), .A1 (n_0_0_283), .A2 (n_0_0_282));
INV_X1 i_0_0_472 (.ZN (n_0_0_280), .A (n_0_0_281));
AOI21_X1 i_0_0_471 (.ZN (n_0_0_279), .A (n_0_0_296), .B1 (n_0_0_344), .B2 (n_0_0_280));
AOI21_X1 i_0_0_470 (.ZN (n_0_0_278), .A (n_0_0_297), .B1 (sps__n7), .B2 (n_0_0_279));
OAI22_X1 i_0_0_469 (.ZN (n_0_148), .A1 (n_0_0_356), .A2 (n_0_0_278), .B1 (sps__n11), .B2 (n_0_0_290));
AOI22_X1 i_0_0_468 (.ZN (n_0_0_277), .A1 (op1[27]), .A2 (spc__n22), .B1 (op1[26]), .B2 (sps__n4));
AOI22_X1 i_0_0_467 (.ZN (n_0_0_276), .A1 (\OP1_complement[27] ), .A2 (spc__n19), .B1 (\OP1_complement[26] ), .B2 (sps__n16));
NAND2_X1 i_0_0_466 (.ZN (n_0_0_275), .A1 (n_0_0_277), .A2 (n_0_0_276));
INV_X1 i_0_0_465 (.ZN (n_0_0_274), .A (n_0_0_275));
AOI21_X1 i_0_0_464 (.ZN (n_0_0_273), .A (n_0_0_296), .B1 (n_0_0_344), .B2 (n_0_0_274));
AOI21_X1 i_0_0_463 (.ZN (n_0_0_272), .A (n_0_0_297), .B1 (sps__n7), .B2 (n_0_0_273));
OAI22_X1 i_0_0_462 (.ZN (n_0_147), .A1 (n_0_0_356), .A2 (n_0_0_272), .B1 (sps__n11), .B2 (n_0_0_284));
AOI22_X1 i_0_0_461 (.ZN (n_0_0_271), .A1 (op1[26]), .A2 (spc__n22), .B1 (op1[25]), .B2 (sps__n4));
AOI22_X1 i_0_0_460 (.ZN (n_0_0_270), .A1 (\OP1_complement[26] ), .A2 (spc__n19), .B1 (\OP1_complement[25] ), .B2 (sps__n16));
NAND2_X1 i_0_0_459 (.ZN (n_0_0_269), .A1 (n_0_0_271), .A2 (n_0_0_270));
INV_X1 i_0_0_458 (.ZN (n_0_0_268), .A (n_0_0_269));
AOI21_X1 i_0_0_457 (.ZN (n_0_0_267), .A (n_0_0_296), .B1 (n_0_0_344), .B2 (n_0_0_268));
AOI22_X1 i_0_0_456 (.ZN (n_0_0_266), .A1 (sps__n1), .A2 (n_0_0_291), .B1 (sps__n7), .B2 (n_0_0_267));
OAI22_X1 i_0_0_455 (.ZN (n_0_146), .A1 (n_0_0_356), .A2 (n_0_0_266), .B1 (sps__n11), .B2 (n_0_0_278));
AOI22_X1 i_0_0_454 (.ZN (n_0_0_265), .A1 (op1[25]), .A2 (spc__n22), .B1 (\OP1_complement[24] ), .B2 (sps__n16));
AOI22_X1 i_0_0_453 (.ZN (n_0_0_264), .A1 (\OP1_complement[25] ), .A2 (spc__n19), .B1 (op1[24]), .B2 (sps__n4));
NAND2_X1 i_0_0_452 (.ZN (n_0_0_263), .A1 (n_0_0_265), .A2 (n_0_0_264));
INV_X1 i_0_0_451 (.ZN (n_0_0_262), .A (n_0_0_263));
AOI21_X1 i_0_0_450 (.ZN (n_0_0_261), .A (n_0_0_296), .B1 (n_0_0_344), .B2 (n_0_0_262));
AOI22_X1 i_0_0_449 (.ZN (n_0_0_260), .A1 (sps__n1), .A2 (n_0_0_285), .B1 (sps__n7), .B2 (n_0_0_261));
OAI22_X1 i_0_0_448 (.ZN (n_0_145), .A1 (n_0_0_356), .A2 (n_0_0_260), .B1 (sps__n11), .B2 (n_0_0_272));
AOI22_X1 i_0_0_447 (.ZN (n_0_0_259), .A1 (op1[24]), .A2 (spc__n22), .B1 (\OP1_complement[24] ), .B2 (spc__n19));
INV_X1 i_0_0_446 (.ZN (n_0_0_258), .A (n_0_0_259));
AOI221_X1 i_0_0_445 (.ZN (n_0_0_257), .A (n_0_0_258), .B1 (op1[23]), .B2 (sps__n4)
    , .C1 (\OP1_complement[23] ), .C2 (sps__n16));
AOI21_X1 i_0_0_444 (.ZN (n_0_0_256), .A (n_0_0_296), .B1 (n_0_0_344), .B2 (n_0_0_257));
AOI22_X1 i_0_0_443 (.ZN (n_0_0_255), .A1 (sps__n7), .A2 (n_0_0_256), .B1 (sps__n1), .B2 (n_0_0_279));
OAI22_X1 i_0_0_442 (.ZN (n_0_144), .A1 (n_0_0_356), .A2 (n_0_0_255), .B1 (sps__n11), .B2 (n_0_0_266));
AOI22_X1 i_0_0_441 (.ZN (n_0_0_254), .A1 (op1[23]), .A2 (spc__n22), .B1 (op1[22]), .B2 (sps__n4));
AOI22_X1 i_0_0_440 (.ZN (n_0_0_253), .A1 (\OP1_complement[23] ), .A2 (spc__n19), .B1 (\OP1_complement[22] ), .B2 (sps__n16));
NAND2_X1 i_0_0_439 (.ZN (n_0_0_252), .A1 (n_0_0_254), .A2 (n_0_0_253));
INV_X1 i_0_0_438 (.ZN (n_0_0_251), .A (n_0_0_252));
AOI21_X1 i_0_0_437 (.ZN (n_0_0_250), .A (n_0_0_296), .B1 (n_0_0_344), .B2 (n_0_0_251));
AOI22_X1 i_0_0_436 (.ZN (n_0_0_249), .A1 (sps__n1), .A2 (n_0_0_273), .B1 (sps__n7), .B2 (n_0_0_250));
OAI22_X1 i_0_0_435 (.ZN (n_0_143), .A1 (n_0_0_356), .A2 (n_0_0_249), .B1 (sps__n11), .B2 (n_0_0_260));
AOI22_X1 i_0_0_434 (.ZN (n_0_0_248), .A1 (op1[22]), .A2 (spc__n22), .B1 (\OP1_complement[21] ), .B2 (sps__n16));
AOI22_X1 i_0_0_433 (.ZN (n_0_0_247), .A1 (\OP1_complement[22] ), .A2 (spc__n19), .B1 (op1[21]), .B2 (sps__n4));
NAND2_X1 i_0_0_432 (.ZN (n_0_0_246), .A1 (n_0_0_248), .A2 (n_0_0_247));
INV_X1 i_0_0_431 (.ZN (n_0_0_245), .A (n_0_0_246));
NOR2_X1 i_0_0_430 (.ZN (n_0_0_244), .A1 (\n[3] ), .A2 (n_0_0_299));
AOI21_X1 i_0_0_429 (.ZN (n_0_0_243), .A (n_0_0_244), .B1 (n_0_0_342), .B2 (n_0_0_293));
OAI21_X1 i_0_0_428 (.ZN (n_0_0_242), .A (n_0_0_243), .B1 (n_0_0_345), .B2 (n_0_0_245));
AOI22_X1 i_0_0_427 (.ZN (n_0_0_241), .A1 (sps__n7), .A2 (n_0_0_242), .B1 (sps__n1), .B2 (n_0_0_267));
OAI22_X1 i_0_0_426 (.ZN (n_0_142), .A1 (n_0_0_356), .A2 (n_0_0_241), .B1 (sps__n11), .B2 (n_0_0_255));
AOI22_X1 i_0_0_425 (.ZN (n_0_0_240), .A1 (op1[21]), .A2 (spc__n22), .B1 (\OP1_complement[20] ), .B2 (sps__n16));
AOI22_X1 i_0_0_424 (.ZN (n_0_0_239), .A1 (\OP1_complement[21] ), .A2 (spc__n19), .B1 (op1[20]), .B2 (sps__n4));
NAND2_X1 i_0_0_423 (.ZN (n_0_0_238), .A1 (n_0_0_240), .A2 (n_0_0_239));
AOI21_X1 i_0_0_422 (.ZN (n_0_0_237), .A (n_0_0_244), .B1 (n_0_0_344), .B2 (n_0_0_238));
OAI21_X1 i_0_0_421 (.ZN (n_0_0_236), .A (n_0_0_237), .B1 (n_0_0_343), .B2 (n_0_0_286));
AOI22_X1 i_0_0_420 (.ZN (n_0_0_235), .A1 (sps__n7), .A2 (n_0_0_236), .B1 (sps__n1), .B2 (n_0_0_261));
OAI22_X1 i_0_0_419 (.ZN (n_0_141), .A1 (n_0_0_356), .A2 (n_0_0_235), .B1 (sps__n11), .B2 (n_0_0_249));
AOI22_X1 i_0_0_418 (.ZN (n_0_0_234), .A1 (\OP1_complement[20] ), .A2 (spc__n19), .B1 (\OP1_complement[19] ), .B2 (sps__n16));
AOI22_X1 i_0_0_417 (.ZN (n_0_0_233), .A1 (op1[20]), .A2 (spc__n22), .B1 (op1[19]), .B2 (sps__n4));
NAND2_X1 i_0_0_416 (.ZN (n_0_0_232), .A1 (n_0_0_234), .A2 (n_0_0_233));
INV_X1 i_0_0_415 (.ZN (n_0_0_231), .A (n_0_0_232));
AOI21_X1 i_0_0_414 (.ZN (n_0_0_230), .A (n_0_0_244), .B1 (n_0_0_342), .B2 (n_0_0_281));
OAI21_X1 i_0_0_413 (.ZN (n_0_0_229), .A (n_0_0_230), .B1 (n_0_0_345), .B2 (n_0_0_231));
AOI22_X1 i_0_0_412 (.ZN (n_0_0_228), .A1 (sps__n7), .A2 (n_0_0_229), .B1 (sps__n1), .B2 (n_0_0_256));
OAI22_X1 i_0_0_411 (.ZN (n_0_140), .A1 (n_0_0_356), .A2 (n_0_0_228), .B1 (sps__n11), .B2 (n_0_0_241));
AOI22_X1 i_0_0_410 (.ZN (n_0_0_227), .A1 (op1[19]), .A2 (spc__n22), .B1 (\OP1_complement[18] ), .B2 (sps__n16));
AOI22_X1 i_0_0_409 (.ZN (n_0_0_226), .A1 (\OP1_complement[19] ), .A2 (spc__n19), .B1 (op1[18]), .B2 (sps__n4));
NAND2_X1 i_0_0_408 (.ZN (n_0_0_225), .A1 (n_0_0_227), .A2 (n_0_0_226));
INV_X1 i_0_0_407 (.ZN (n_0_0_224), .A (n_0_0_225));
AOI21_X1 i_0_0_406 (.ZN (n_0_0_223), .A (n_0_0_244), .B1 (n_0_0_342), .B2 (n_0_0_275));
OAI21_X1 i_0_0_405 (.ZN (n_0_0_222), .A (n_0_0_223), .B1 (n_0_0_345), .B2 (n_0_0_224));
AOI22_X1 i_0_0_404 (.ZN (n_0_0_221), .A1 (sps__n7), .A2 (n_0_0_222), .B1 (sps__n1), .B2 (n_0_0_250));
OAI22_X1 i_0_0_403 (.ZN (n_0_139), .A1 (n_0_0_356), .A2 (n_0_0_221), .B1 (sps__n11), .B2 (n_0_0_235));
AOI22_X1 i_0_0_402 (.ZN (n_0_0_220), .A1 (\OP1_complement[18] ), .A2 (spc__n19), .B1 (\OP1_complement[17] ), .B2 (sps__n16));
AOI22_X1 i_0_0_401 (.ZN (n_0_0_219), .A1 (op1[18]), .A2 (spc__n22), .B1 (op1[17]), .B2 (sps__n4));
NAND2_X1 i_0_0_400 (.ZN (n_0_0_218), .A1 (n_0_0_220), .A2 (n_0_0_219));
INV_X1 i_0_0_399 (.ZN (n_0_0_217), .A (n_0_0_218));
AOI21_X1 i_0_0_398 (.ZN (n_0_0_216), .A (n_0_0_244), .B1 (n_0_0_342), .B2 (n_0_0_269));
OAI21_X1 i_0_0_397 (.ZN (n_0_0_215), .A (n_0_0_216), .B1 (n_0_0_345), .B2 (n_0_0_217));
AOI22_X1 i_0_0_396 (.ZN (n_0_0_214), .A1 (sps__n1), .A2 (n_0_0_242), .B1 (sps__n7), .B2 (n_0_0_215));
OAI22_X1 i_0_0_395 (.ZN (n_0_138), .A1 (n_0_0_356), .A2 (n_0_0_214), .B1 (sps__n11), .B2 (n_0_0_228));
AOI22_X1 i_0_0_394 (.ZN (n_0_0_213), .A1 (op1[17]), .A2 (spc__n22), .B1 (op1[16]), .B2 (sps__n4));
AOI22_X1 i_0_0_393 (.ZN (n_0_0_212), .A1 (\OP1_complement[17] ), .A2 (spc__n19), .B1 (\OP1_complement[16] ), .B2 (sps__n16));
NAND2_X1 i_0_0_392 (.ZN (n_0_0_211), .A1 (n_0_0_213), .A2 (n_0_0_212));
INV_X1 i_0_0_391 (.ZN (n_0_0_210), .A (n_0_0_211));
AOI21_X1 i_0_0_390 (.ZN (n_0_0_209), .A (n_0_0_244), .B1 (n_0_0_342), .B2 (n_0_0_263));
OAI21_X1 i_0_0_389 (.ZN (n_0_0_208), .A (n_0_0_209), .B1 (n_0_0_345), .B2 (n_0_0_210));
AOI22_X1 i_0_0_388 (.ZN (n_0_0_207), .A1 (sps__n7), .A2 (n_0_0_208), .B1 (sps__n1), .B2 (n_0_0_236));
OAI22_X1 i_0_0_387 (.ZN (n_0_137), .A1 (n_0_0_356), .A2 (n_0_0_207), .B1 (sps__n11), .B2 (n_0_0_221));
AOI22_X1 i_0_0_386 (.ZN (n_0_0_206), .A1 (\OP1_complement[16] ), .A2 (spc__n19), .B1 (\OP1_complement[15] ), .B2 (sps__n16));
AOI22_X1 i_0_0_385 (.ZN (n_0_0_205), .A1 (op1[16]), .A2 (spc__n22), .B1 (op1[15]), .B2 (sps__n4));
NAND2_X1 i_0_0_384 (.ZN (n_0_0_204), .A1 (n_0_0_206), .A2 (n_0_0_205));
AOI21_X1 i_0_0_383 (.ZN (n_0_0_203), .A (n_0_0_244), .B1 (n_0_0_344), .B2 (n_0_0_204));
OAI21_X1 i_0_0_382 (.ZN (n_0_0_202), .A (n_0_0_203), .B1 (n_0_0_343), .B2 (n_0_0_257));
AOI22_X1 i_0_0_381 (.ZN (n_0_0_201), .A1 (sps__n1), .A2 (n_0_0_229), .B1 (sps__n7), .B2 (n_0_0_202));
OAI22_X1 i_0_0_380 (.ZN (n_0_136), .A1 (n_0_0_356), .A2 (n_0_0_201), .B1 (sps__n11), .B2 (n_0_0_214));
AOI22_X1 i_0_0_379 (.ZN (n_0_0_200), .A1 (\OP1_complement[15] ), .A2 (spc__n19), .B1 (\OP1_complement[14] ), .B2 (sps__n16));
AOI22_X1 i_0_0_378 (.ZN (n_0_0_199), .A1 (op1[15]), .A2 (spc__n22), .B1 (op1[14]), .B2 (sps__n4));
NAND2_X1 i_0_0_377 (.ZN (n_0_0_198), .A1 (n_0_0_200), .A2 (n_0_0_199));
AOI21_X1 i_0_0_376 (.ZN (n_0_0_197), .A (n_0_0_244), .B1 (n_0_0_344), .B2 (n_0_0_198));
OAI21_X1 i_0_0_375 (.ZN (n_0_0_196), .A (n_0_0_197), .B1 (n_0_0_343), .B2 (n_0_0_251));
AOI22_X1 i_0_0_374 (.ZN (n_0_0_195), .A1 (sps__n1), .A2 (n_0_0_222), .B1 (sps__n7), .B2 (n_0_0_196));
OAI22_X1 i_0_0_373 (.ZN (n_0_135), .A1 (n_0_0_356), .A2 (n_0_0_195), .B1 (sps__n11), .B2 (n_0_0_207));
NOR2_X1 i_0_0_372 (.ZN (n_0_0_194), .A1 (n_0_0_340), .A2 (n_0_89));
AOI22_X1 i_0_0_371 (.ZN (n_0_0_193), .A1 (\OP1_complement[14] ), .A2 (spc__n19), .B1 (\OP1_complement[13] ), .B2 (sps__n16));
AOI22_X1 i_0_0_370 (.ZN (n_0_0_192), .A1 (op1[14]), .A2 (spc__n22), .B1 (op1[13]), .B2 (sps__n4));
NAND2_X1 i_0_0_369 (.ZN (n_0_0_191), .A1 (n_0_0_193), .A2 (n_0_0_192));
OAI22_X1 i_0_0_368 (.ZN (n_0_0_190), .A1 (n_0_0_343), .A2 (n_0_0_246), .B1 (n_0_0_345), .B2 (n_0_0_191));
AOI211_X1 i_0_0_367 (.ZN (n_0_0_189), .A (n_0_0_194), .B (n_0_0_190), .C1 (n_0_0_349), .C2 (n_0_0_292));
AOI22_X1 i_0_0_366 (.ZN (n_0_0_188), .A1 (sps__n7), .A2 (n_0_0_189), .B1 (sps__n1), .B2 (n_0_0_215));
OAI22_X1 i_0_0_365 (.ZN (n_0_134), .A1 (sps__n11), .A2 (n_0_0_201), .B1 (n_0_0_356), .B2 (n_0_0_188));
AOI22_X1 i_0_0_364 (.ZN (n_0_0_187), .A1 (\OP1_complement[13] ), .A2 (spc__n19), .B1 (\OP1_complement[12] ), .B2 (sps__n16));
AOI22_X1 i_0_0_363 (.ZN (n_0_0_186), .A1 (op1[13]), .A2 (spc__n22), .B1 (op1[12]), .B2 (sps__n4));
NAND2_X1 i_0_0_362 (.ZN (n_0_0_185), .A1 (n_0_0_187), .A2 (n_0_0_186));
INV_X1 i_0_0_361 (.ZN (n_0_0_184), .A (n_0_0_185));
OAI22_X1 i_0_0_360 (.ZN (n_0_0_183), .A1 (n_0_0_350), .A2 (n_0_0_287), .B1 (n_0_0_343), .B2 (n_0_0_238));
AOI211_X1 i_0_0_359 (.ZN (n_0_0_182), .A (n_0_0_194), .B (n_0_0_183), .C1 (n_0_0_344), .C2 (n_0_0_184));
AOI22_X1 i_0_0_358 (.ZN (n_0_0_181), .A1 (sps__n7), .A2 (n_0_0_182), .B1 (sps__n1), .B2 (n_0_0_208));
OAI22_X1 i_0_0_357 (.ZN (n_0_133), .A1 (n_0_0_356), .A2 (n_0_0_181), .B1 (sps__n11), .B2 (n_0_0_195));
AOI22_X1 i_0_0_356 (.ZN (n_0_0_180), .A1 (op1[12]), .A2 (spc__n22), .B1 (\OP1_complement[11] ), .B2 (sps__n16));
AOI22_X1 i_0_0_355 (.ZN (n_0_0_179), .A1 (\OP1_complement[12] ), .A2 (spc__n19), .B1 (op1[11]), .B2 (sps__n4));
NAND2_X1 i_0_0_354 (.ZN (n_0_0_178), .A1 (n_0_0_180), .A2 (n_0_0_179));
INV_X1 i_0_0_353 (.ZN (n_0_0_177), .A (n_0_0_178));
OAI22_X1 i_0_0_352 (.ZN (n_0_0_176), .A1 (n_0_0_343), .A2 (n_0_0_232), .B1 (n_0_0_345), .B2 (n_0_0_178));
AOI211_X1 i_0_0_351 (.ZN (n_0_0_175), .A (n_0_0_194), .B (n_0_0_176), .C1 (n_0_0_349), .C2 (n_0_0_280));
AOI22_X1 i_0_0_350 (.ZN (n_0_0_174), .A1 (sps__n7), .A2 (n_0_0_175), .B1 (sps__n1), .B2 (n_0_0_202));
OAI22_X1 i_0_0_349 (.ZN (n_0_132), .A1 (n_0_0_356), .A2 (n_0_0_174), .B1 (sps__n11), .B2 (n_0_0_188));
AOI22_X1 i_0_0_348 (.ZN (n_0_0_173), .A1 (\OP1_complement[11] ), .A2 (spc__n19), .B1 (\OP1_complement[10] ), .B2 (sps__n16));
AOI22_X1 i_0_0_347 (.ZN (n_0_0_172), .A1 (op1[11]), .A2 (spc__n22), .B1 (op1[10]), .B2 (sps__n4));
NAND2_X1 i_0_0_346 (.ZN (n_0_0_171), .A1 (n_0_0_173), .A2 (n_0_0_172));
INV_X1 i_0_0_345 (.ZN (n_0_0_170), .A (n_0_0_171));
OAI22_X1 i_0_0_344 (.ZN (n_0_0_169), .A1 (n_0_0_350), .A2 (n_0_0_275), .B1 (n_0_0_343), .B2 (n_0_0_225));
AOI211_X1 i_0_0_343 (.ZN (n_0_0_168), .A (n_0_0_194), .B (n_0_0_169), .C1 (n_0_0_344), .C2 (n_0_0_170));
AOI22_X1 i_0_0_342 (.ZN (n_0_0_167), .A1 (sps__n7), .A2 (n_0_0_168), .B1 (sps__n1), .B2 (n_0_0_196));
OAI22_X1 i_0_0_341 (.ZN (n_0_131), .A1 (n_0_0_356), .A2 (n_0_0_167), .B1 (sps__n11), .B2 (n_0_0_181));
AOI22_X1 i_0_0_340 (.ZN (n_0_0_166), .A1 (\OP1_complement[10] ), .A2 (spc__n19), .B1 (\OP1_complement[9] ), .B2 (sps__n16));
AOI22_X1 i_0_0_339 (.ZN (n_0_0_165), .A1 (op1[10]), .A2 (spc__n22), .B1 (op1[9]), .B2 (sps__n4));
NAND2_X1 i_0_0_338 (.ZN (n_0_0_164), .A1 (n_0_0_166), .A2 (n_0_0_165));
OAI22_X1 i_0_0_337 (.ZN (n_0_0_163), .A1 (n_0_0_343), .A2 (n_0_0_218), .B1 (n_0_0_345), .B2 (n_0_0_164));
AOI211_X1 i_0_0_336 (.ZN (n_0_0_162), .A (n_0_0_194), .B (n_0_0_163), .C1 (n_0_0_349), .C2 (n_0_0_268));
AOI22_X1 i_0_0_335 (.ZN (n_0_0_161), .A1 (sps__n1), .A2 (n_0_0_189), .B1 (sps__n7), .B2 (n_0_0_162));
OAI22_X1 i_0_0_334 (.ZN (n_0_130), .A1 (sps__n11), .A2 (n_0_0_174), .B1 (n_0_0_356), .B2 (n_0_0_161));
AOI22_X1 i_0_0_333 (.ZN (n_0_0_160), .A1 (\OP1_complement[9] ), .A2 (spc__n19), .B1 (\OP1_complement[8] ), .B2 (sps__n16));
AOI22_X1 i_0_0_332 (.ZN (n_0_0_159), .A1 (op1[9]), .A2 (spc__n22), .B1 (op1[8]), .B2 (sps__n4));
NAND2_X1 i_0_0_331 (.ZN (n_0_0_158), .A1 (n_0_0_160), .A2 (n_0_0_159));
INV_X1 i_0_0_330 (.ZN (n_0_0_157), .A (n_0_0_158));
OAI22_X1 i_0_0_329 (.ZN (n_0_0_156), .A1 (n_0_0_343), .A2 (n_0_0_211), .B1 (n_0_0_350), .B2 (n_0_0_263));
AOI211_X1 i_0_0_328 (.ZN (n_0_0_155), .A (n_0_0_194), .B (n_0_0_156), .C1 (n_0_0_344), .C2 (n_0_0_157));
AOI22_X1 i_0_0_327 (.ZN (n_0_0_154), .A1 (sps__n1), .A2 (n_0_0_182), .B1 (sps__n7), .B2 (n_0_0_155));
OAI22_X1 i_0_0_326 (.ZN (n_0_129), .A1 (sps__n11), .A2 (n_0_0_167), .B1 (n_0_0_356), .B2 (n_0_0_154));
AOI22_X1 i_0_0_325 (.ZN (n_0_0_153), .A1 (\OP1_complement[8] ), .A2 (spc__n19), .B1 (\OP1_complement[7] ), .B2 (sps__n16));
AOI22_X1 i_0_0_324 (.ZN (n_0_0_152), .A1 (op1[8]), .A2 (spc__n22), .B1 (op1[7]), .B2 (sps__n4));
NAND2_X1 i_0_0_323 (.ZN (n_0_0_151), .A1 (n_0_0_153), .A2 (n_0_0_152));
INV_X1 i_0_0_322 (.ZN (n_0_0_150), .A (n_0_0_151));
AOI22_X1 i_0_0_321 (.ZN (n_0_0_149), .A1 (n_0_0_359), .A2 (n_0_0_257), .B1 (\n[3] ), .B2 (n_0_0_150));
AOI22_X1 i_0_0_320 (.ZN (n_0_0_148), .A1 (\n[2] ), .A2 (n_0_0_149), .B1 (n_0_0_342), .B2 (n_0_0_204));
OAI21_X1 i_0_0_319 (.ZN (n_0_0_147), .A (n_0_0_148), .B1 (n_0_0_340), .B2 (n_0_0_299));
AOI22_X1 i_0_0_318 (.ZN (n_0_0_146), .A1 (sps__n1), .A2 (n_0_0_175), .B1 (sps__n7), .B2 (n_0_0_147));
OAI22_X1 i_0_0_317 (.ZN (n_0_128), .A1 (sps__n10), .A2 (n_0_0_161), .B1 (n_0_0_356), .B2 (n_0_0_146));
AOI22_X1 i_0_0_316 (.ZN (n_0_0_145), .A1 (op1[6]), .A2 (sps__n4), .B1 (\OP1_complement[6] ), .B2 (sps__n16));
AOI22_X1 i_0_0_315 (.ZN (n_0_0_144), .A1 (op1[7]), .A2 (spc__n22), .B1 (\OP1_complement[7] ), .B2 (spc__n19));
NAND2_X1 i_0_0_314 (.ZN (n_0_0_143), .A1 (n_0_0_145), .A2 (n_0_0_144));
OAI22_X1 i_0_0_313 (.ZN (n_0_0_142), .A1 (n_0_0_358), .A2 (n_0_0_143), .B1 (\n[2] ), .B2 (n_0_0_198));
INV_X1 i_0_0_312 (.ZN (n_0_0_141), .A (n_0_0_142));
AOI221_X1 i_0_0_311 (.ZN (n_0_0_140), .A (n_0_0_194), .B1 (n_0_0_349), .B2 (n_0_0_251)
    , .C1 (\n[3] ), .C2 (n_0_0_142));
AOI22_X1 i_0_0_310 (.ZN (n_0_0_139), .A1 (sps__n1), .A2 (n_0_0_168), .B1 (sps__n7), .B2 (n_0_0_140));
OAI22_X1 i_0_0_309 (.ZN (n_0_127), .A1 (n_0_0_356), .A2 (n_0_0_139), .B1 (sps__n10), .B2 (n_0_0_154));
AOI22_X1 i_0_0_308 (.ZN (n_0_0_138), .A1 (op1[5]), .A2 (sps__n4), .B1 (\OP1_complement[5] ), .B2 (sps__n16));
AOI22_X1 i_0_0_307 (.ZN (n_0_0_137), .A1 (op1[6]), .A2 (spc__n22), .B1 (\OP1_complement[6] ), .B2 (spc__n19));
NAND2_X1 i_0_0_306 (.ZN (n_0_0_136), .A1 (n_0_0_138), .A2 (n_0_0_137));
OAI22_X1 i_0_0_305 (.ZN (n_0_0_135), .A1 (n_0_0_358), .A2 (n_0_0_136), .B1 (\n[2] ), .B2 (n_0_0_191));
INV_X1 i_0_0_304 (.ZN (n_0_0_134), .A (n_0_0_135));
AOI222_X1 i_0_0_303 (.ZN (n_0_0_133), .A1 (n_0_0_339), .A2 (n_0_0_292), .B1 (n_0_0_349)
    , .B2 (n_0_0_245), .C1 (\n[3] ), .C2 (n_0_0_135));
AOI22_X1 i_0_0_302 (.ZN (n_0_0_132), .A1 (sps__n7), .A2 (n_0_0_133), .B1 (sps__n1), .B2 (n_0_0_162));
OAI22_X1 i_0_0_301 (.ZN (n_0_126), .A1 (n_0_0_356), .A2 (n_0_0_132), .B1 (sps__n10), .B2 (n_0_0_146));
AOI22_X1 i_0_0_300 (.ZN (n_0_0_131), .A1 (\OP1_complement[5] ), .A2 (spc__n19), .B1 (\OP1_complement[4] ), .B2 (sps__n16));
AOI22_X1 i_0_0_299 (.ZN (n_0_0_130), .A1 (op1[5]), .A2 (spc__n22), .B1 (op1[4]), .B2 (sps__n4));
NAND2_X1 i_0_0_298 (.ZN (n_0_0_129), .A1 (n_0_0_131), .A2 (n_0_0_130));
NOR2_X1 i_0_0_297 (.ZN (n_0_0_128), .A1 (n_0_0_358), .A2 (n_0_0_129));
AOI21_X1 i_0_0_296 (.ZN (n_0_0_127), .A (n_0_0_128), .B1 (n_0_0_358), .B2 (n_0_0_184));
OAI222_X1 i_0_0_295 (.ZN (n_0_0_126), .A1 (n_0_0_340), .A2 (n_0_0_287), .B1 (n_0_0_350)
    , .B2 (n_0_0_238), .C1 (n_0_0_359), .C2 (n_0_0_127));
NAND2_X1 i_0_0_294 (.ZN (n_0_0_125), .A1 (sps__n1), .A2 (n_0_0_155));
OAI21_X1 i_0_0_293 (.ZN (n_0_0_124), .A (n_0_0_125), .B1 (sps__n1), .B2 (n_0_0_126));
NAND2_X1 i_0_0_292 (.ZN (n_0_0_123), .A1 (sps__n10), .A2 (n_0_0_124));
OAI21_X1 i_0_0_291 (.ZN (n_0_125), .A (n_0_0_123), .B1 (sps__n10), .B2 (n_0_0_139));
AOI22_X1 i_0_0_290 (.ZN (n_0_0_122), .A1 (op1[3]), .A2 (sps__n4), .B1 (\OP1_complement[3] ), .B2 (sps__n16));
AOI22_X1 i_0_0_289 (.ZN (n_0_0_121), .A1 (op1[4]), .A2 (spc__n22), .B1 (\OP1_complement[4] ), .B2 (spc__n19));
NAND2_X1 i_0_0_288 (.ZN (n_0_0_120), .A1 (n_0_0_122), .A2 (n_0_0_121));
INV_X1 i_0_0_287 (.ZN (n_0_0_119), .A (n_0_0_120));
AOI22_X1 i_0_0_286 (.ZN (n_0_0_118), .A1 (n_0_0_359), .A2 (n_0_0_231), .B1 (\n[3] ), .B2 (n_0_0_119));
INV_X1 i_0_0_285 (.ZN (n_0_0_117), .A (n_0_0_118));
AOI222_X1 i_0_0_284 (.ZN (n_0_0_116), .A1 (n_0_0_339), .A2 (n_0_0_280), .B1 (n_0_0_342)
    , .B2 (n_0_0_177), .C1 (\n[2] ), .C2 (n_0_0_117));
AOI22_X1 i_0_0_283 (.ZN (n_0_0_115), .A1 (sps__n7), .A2 (n_0_0_116), .B1 (sps__n1), .B2 (n_0_0_147));
OAI22_X1 i_0_0_282 (.ZN (n_0_124), .A1 (n_0_0_356), .A2 (n_0_0_115), .B1 (sps__n10), .B2 (n_0_0_132));
AOI22_X1 i_0_0_281 (.ZN (n_0_0_114), .A1 (\OP1_complement[3] ), .A2 (spc__n19), .B1 (\OP1_complement[2] ), .B2 (sps__n16));
AOI22_X1 i_0_0_280 (.ZN (n_0_0_113), .A1 (op1[3]), .A2 (spc__n22), .B1 (op1[2]), .B2 (sps__n4));
NAND2_X1 i_0_0_279 (.ZN (n_0_0_112), .A1 (n_0_0_114), .A2 (n_0_0_113));
NOR2_X1 i_0_0_278 (.ZN (n_0_0_111), .A1 (n_0_0_358), .A2 (n_0_0_112));
AOI21_X1 i_0_0_277 (.ZN (n_0_0_110), .A (n_0_0_111), .B1 (n_0_0_358), .B2 (n_0_0_170));
OAI222_X1 i_0_0_276 (.ZN (n_0_0_109), .A1 (n_0_0_350), .A2 (n_0_0_225), .B1 (n_0_0_340)
    , .B2 (n_0_0_275), .C1 (n_0_0_359), .C2 (n_0_0_110));
NAND2_X1 i_0_0_275 (.ZN (n_0_0_108), .A1 (sps__n1), .A2 (n_0_0_140));
OAI21_X1 i_0_0_274 (.ZN (n_0_0_107), .A (n_0_0_108), .B1 (sps__n1), .B2 (n_0_0_109));
AOI22_X1 i_0_0_273 (.ZN (n_0_0_106), .A1 (n_0_0_356), .A2 (n_0_0_124), .B1 (sps__n10), .B2 (n_0_0_107));
INV_X1 i_0_0_272 (.ZN (n_0_123), .A (n_0_0_106));
AOI22_X1 i_0_0_271 (.ZN (n_0_0_105), .A1 (\OP1_complement[2] ), .A2 (spc__n19), .B1 (\OP1_complement[1] ), .B2 (sps__n16));
AOI22_X1 i_0_0_270 (.ZN (n_0_0_104), .A1 (op1[2]), .A2 (spc__n22), .B1 (op1[1]), .B2 (sps__n4));
NAND2_X1 i_0_0_269 (.ZN (n_0_0_103), .A1 (n_0_0_105), .A2 (n_0_0_104));
OAI22_X1 i_0_0_268 (.ZN (n_0_0_102), .A1 (n_0_0_358), .A2 (n_0_0_103), .B1 (\n[2] ), .B2 (n_0_0_164));
INV_X1 i_0_0_267 (.ZN (n_0_0_101), .A (n_0_0_102));
AOI222_X1 i_0_0_266 (.ZN (n_0_0_100), .A1 (n_0_0_339), .A2 (n_0_0_268), .B1 (n_0_0_349)
    , .B2 (n_0_0_217), .C1 (\n[3] ), .C2 (n_0_0_102));
AOI22_X1 i_0_0_265 (.ZN (n_0_0_99), .A1 (sps__n7), .A2 (n_0_0_100), .B1 (sps__n1), .B2 (n_0_0_133));
OAI22_X1 i_0_0_264 (.ZN (n_0_122), .A1 (sps__n10), .A2 (n_0_0_115), .B1 (n_0_0_356), .B2 (n_0_0_99));
AOI22_X1 i_0_0_263 (.ZN (n_0_0_98), .A1 (\OP1_complement[1] ), .A2 (spc__n19), .B1 (\OP1_complement[0] ), .B2 (sps__n16));
AOI22_X1 i_0_0_262 (.ZN (n_0_0_97), .A1 (op1[1]), .A2 (spc__n22), .B1 (op1[0]), .B2 (sps__n4));
NAND2_X1 i_0_0_261 (.ZN (n_0_0_96), .A1 (n_0_0_98), .A2 (n_0_0_97));
NOR2_X1 i_0_0_260 (.ZN (n_0_0_95), .A1 (n_0_0_358), .A2 (n_0_0_96));
AOI21_X1 i_0_0_259 (.ZN (n_0_0_94), .A (n_0_0_95), .B1 (n_0_0_358), .B2 (n_0_0_157));
OAI222_X1 i_0_0_258 (.ZN (n_0_0_93), .A1 (n_0_0_340), .A2 (n_0_0_263), .B1 (n_0_0_350)
    , .B2 (n_0_0_211), .C1 (n_0_0_359), .C2 (n_0_0_94));
AOI22_X1 i_0_0_257 (.ZN (n_0_0_92), .A1 (sps__n1), .A2 (n_0_0_126), .B1 (sps__n7), .B2 (n_0_0_93));
AOI22_X1 i_0_0_256 (.ZN (n_0_0_91), .A1 (sps__n10), .A2 (n_0_0_92), .B1 (n_0_0_356), .B2 (n_0_0_107));
INV_X1 i_0_0_255 (.ZN (n_0_121), .A (n_0_0_91));
AOI22_X1 i_0_0_254 (.ZN (n_0_0_90), .A1 (\OP1_complement[0] ), .A2 (spc__n19), .B1 (op1[0]), .B2 (spc__n22));
INV_X1 i_0_0_253 (.ZN (n_0_0_89), .A (n_0_0_90));
NAND2_X1 i_0_0_252 (.ZN (n_0_0_88), .A1 (n_0_0_359), .A2 (n_0_0_204));
OAI21_X1 i_0_0_251 (.ZN (n_0_0_87), .A (n_0_0_88), .B1 (n_0_0_359), .B2 (n_0_0_90));
AOI22_X1 i_0_0_250 (.ZN (n_0_0_86), .A1 (\n[2] ), .A2 (n_0_0_87), .B1 (n_0_0_358), .B2 (n_0_0_149));
NAND2_X1 i_0_0_249 (.ZN (n_0_0_85), .A1 (sps__n1), .A2 (n_0_0_116));
OAI21_X1 i_0_0_248 (.ZN (n_0_0_84), .A (n_0_0_85), .B1 (sps__n1), .B2 (n_0_0_86));
NAND2_X1 i_0_0_247 (.ZN (n_0_0_83), .A1 (sps__n10), .A2 (n_0_0_84));
OAI21_X1 i_0_0_246 (.ZN (n_0_120), .A (n_0_0_83), .B1 (sps__n10), .B2 (n_0_0_99));
AOI222_X1 i_0_0_245 (.ZN (n_0_0_82), .A1 (n_0_0_339), .A2 (n_0_0_252), .B1 (n_0_0_342)
    , .B2 (n_0_0_143), .C1 (n_0_0_349), .C2 (n_0_0_198));
AOI22_X1 i_0_0_244 (.ZN (n_0_0_81), .A1 (sps__n1), .A2 (n_0_0_109), .B1 (sps__n7), .B2 (n_0_0_82));
AOI22_X1 i_0_0_243 (.ZN (n_0_0_80), .A1 (n_0_0_356), .A2 (n_0_0_92), .B1 (sps__n10), .B2 (n_0_0_81));
INV_X1 i_0_0_242 (.ZN (n_0_119), .A (n_0_0_80));
AOI22_X1 i_0_0_241 (.ZN (n_0_0_79), .A1 (n_0_0_342), .A2 (n_0_0_136), .B1 (n_0_0_349), .B2 (n_0_0_191));
OAI21_X1 i_0_0_240 (.ZN (n_0_0_78), .A (n_0_0_79), .B1 (n_0_0_340), .B2 (n_0_0_245));
AOI22_X1 i_0_0_239 (.ZN (n_0_0_77), .A1 (sps__n1), .A2 (n_0_0_100), .B1 (sps__n7), .B2 (n_0_0_78));
NAND2_X1 i_0_0_238 (.ZN (n_0_0_76), .A1 (n_0_0_356), .A2 (n_0_0_84));
OAI21_X1 i_0_0_237 (.ZN (n_0_118), .A (n_0_0_76), .B1 (n_0_0_356), .B2 (n_0_0_77));
AOI222_X1 i_0_0_236 (.ZN (n_0_0_75), .A1 (n_0_0_339), .A2 (n_0_0_238), .B1 (n_0_0_342)
    , .B2 (n_0_0_129), .C1 (n_0_0_349), .C2 (n_0_0_185));
AOI22_X1 i_0_0_235 (.ZN (n_0_0_74), .A1 (sps__n1), .A2 (n_0_0_93), .B1 (sps__n7), .B2 (n_0_0_75));
AOI22_X1 i_0_0_234 (.ZN (n_0_0_73), .A1 (sps__n10), .A2 (n_0_0_74), .B1 (n_0_0_356), .B2 (n_0_0_81));
INV_X1 i_0_0_233 (.ZN (n_0_117), .A (n_0_0_73));
AOI22_X1 i_0_0_232 (.ZN (n_0_0_72), .A1 (n_0_0_358), .A2 (n_0_0_118), .B1 (n_0_0_349), .B2 (n_0_0_178));
OAI22_X1 i_0_0_231 (.ZN (n_0_0_71), .A1 (sps__n1), .A2 (n_0_0_72), .B1 (sps__n7), .B2 (n_0_0_86));
NAND2_X1 i_0_0_230 (.ZN (n_0_0_70), .A1 (sps__n11), .A2 (n_0_0_71));
OAI21_X1 i_0_0_229 (.ZN (n_0_116), .A (n_0_0_70), .B1 (sps__n11), .B2 (n_0_0_77));
AOI22_X1 i_0_0_228 (.ZN (n_0_0_69), .A1 (n_0_0_342), .A2 (n_0_0_112), .B1 (n_0_0_349), .B2 (n_0_0_171));
OAI21_X1 i_0_0_227 (.ZN (n_0_0_68), .A (n_0_0_69), .B1 (n_0_0_340), .B2 (n_0_0_224));
NAND2_X1 i_0_0_226 (.ZN (n_0_0_67), .A1 (sps__n7), .A2 (n_0_0_68));
OAI21_X1 i_0_0_225 (.ZN (n_0_0_66), .A (n_0_0_67), .B1 (sps__n7), .B2 (n_0_0_82));
AOI22_X1 i_0_0_224 (.ZN (n_0_0_65), .A1 (n_0_0_356), .A2 (n_0_0_74), .B1 (sps__n11), .B2 (n_0_0_66));
INV_X1 i_0_0_223 (.ZN (n_0_115), .A (n_0_0_65));
AOI22_X1 i_0_0_222 (.ZN (n_0_0_64), .A1 (n_0_0_349), .A2 (n_0_0_164), .B1 (n_0_0_342), .B2 (n_0_0_103));
OAI21_X1 i_0_0_221 (.ZN (n_0_0_63), .A (n_0_0_64), .B1 (n_0_0_340), .B2 (n_0_0_217));
AOI22_X1 i_0_0_220 (.ZN (n_0_0_62), .A1 (sps__n7), .A2 (n_0_0_63), .B1 (sps__n1), .B2 (n_0_0_78));
NAND2_X1 i_0_0_219 (.ZN (n_0_0_61), .A1 (n_0_0_356), .A2 (n_0_0_71));
OAI21_X1 i_0_0_218 (.ZN (n_0_114), .A (n_0_0_61), .B1 (n_0_0_356), .B2 (n_0_0_62));
AOI22_X1 i_0_0_217 (.ZN (n_0_0_60), .A1 (n_0_0_349), .A2 (n_0_0_158), .B1 (n_0_0_342), .B2 (n_0_0_96));
OAI21_X1 i_0_0_216 (.ZN (n_0_0_59), .A (n_0_0_60), .B1 (n_0_0_340), .B2 (n_0_0_210));
NAND2_X1 i_0_0_215 (.ZN (n_0_0_58), .A1 (sps__n7), .A2 (n_0_0_59));
OAI21_X1 i_0_0_214 (.ZN (n_0_0_57), .A (n_0_0_58), .B1 (sps__n7), .B2 (n_0_0_75));
AOI22_X1 i_0_0_213 (.ZN (n_0_0_56), .A1 (n_0_0_356), .A2 (n_0_0_66), .B1 (sps__n11), .B2 (n_0_0_57));
INV_X1 i_0_0_212 (.ZN (n_0_113), .A (n_0_0_56));
AOI22_X1 i_0_0_211 (.ZN (n_0_0_55), .A1 (n_0_0_358), .A2 (n_0_0_87), .B1 (n_0_0_349), .B2 (n_0_0_151));
AOI22_X1 i_0_0_210 (.ZN (n_0_0_54), .A1 (sps__n1), .A2 (n_0_0_72), .B1 (sps__n7), .B2 (n_0_0_55));
NAND2_X1 i_0_0_209 (.ZN (n_0_0_53), .A1 (sps__n11), .A2 (n_0_0_54));
OAI21_X1 i_0_0_208 (.ZN (n_0_112), .A (n_0_0_53), .B1 (sps__n11), .B2 (n_0_0_62));
NOR2_X1 i_0_0_207 (.ZN (n_0_0_52), .A1 (\n[3] ), .A2 (sps__n1));
AOI22_X1 i_0_0_206 (.ZN (n_0_0_51), .A1 (sps__n1), .A2 (n_0_0_68), .B1 (n_0_0_141), .B2 (n_0_0_52));
NAND2_X1 i_0_0_205 (.ZN (n_0_0_50), .A1 (n_0_0_356), .A2 (n_0_0_57));
OAI21_X1 i_0_0_204 (.ZN (n_0_111), .A (n_0_0_50), .B1 (n_0_0_356), .B2 (n_0_0_51));
AOI22_X1 i_0_0_203 (.ZN (n_0_0_49), .A1 (sps__n1), .A2 (n_0_0_63), .B1 (n_0_0_134), .B2 (n_0_0_52));
NAND2_X1 i_0_0_202 (.ZN (n_0_0_48), .A1 (n_0_0_356), .A2 (n_0_0_54));
OAI21_X1 i_0_0_201 (.ZN (n_0_110), .A (n_0_0_48), .B1 (n_0_0_356), .B2 (n_0_0_49));
AOI22_X1 i_0_0_200 (.ZN (n_0_0_47), .A1 (sps__n1), .A2 (n_0_0_59), .B1 (n_0_0_127), .B2 (n_0_0_52));
OAI22_X1 i_0_0_199 (.ZN (n_0_109), .A1 (sps__n11), .A2 (n_0_0_51), .B1 (n_0_0_356), .B2 (n_0_0_47));
AOI22_X1 i_0_0_198 (.ZN (n_0_0_46), .A1 (\n[2] ), .A2 (n_0_0_119), .B1 (n_0_0_358), .B2 (n_0_0_177));
NAND2_X1 i_0_0_197 (.ZN (n_0_0_45), .A1 (n_0_0_52), .A2 (n_0_0_46));
OAI21_X1 i_0_0_196 (.ZN (n_0_0_44), .A (n_0_0_45), .B1 (sps__n7), .B2 (n_0_0_55));
NAND2_X1 i_0_0_195 (.ZN (n_0_0_43), .A1 (sps__n11), .A2 (n_0_0_44));
OAI21_X1 i_0_0_194 (.ZN (n_0_108), .A (n_0_0_43), .B1 (sps__n11), .B2 (n_0_0_49));
AOI22_X1 i_0_0_193 (.ZN (n_0_0_42), .A1 (n_0_0_110), .A2 (n_0_0_52), .B1 (n_0_0_316), .B2 (n_0_0_141));
OAI22_X1 i_0_0_192 (.ZN (n_0_107), .A1 (sps__n11), .A2 (n_0_0_47), .B1 (n_0_0_356), .B2 (n_0_0_42));
AOI22_X1 i_0_0_191 (.ZN (n_0_0_41), .A1 (n_0_0_101), .A2 (n_0_0_52), .B1 (n_0_0_316), .B2 (n_0_0_134));
NAND2_X1 i_0_0_190 (.ZN (n_0_0_40), .A1 (n_0_0_356), .A2 (n_0_0_44));
OAI21_X1 i_0_0_189 (.ZN (n_0_106), .A (n_0_0_40), .B1 (n_0_0_356), .B2 (n_0_0_41));
AOI22_X1 i_0_0_188 (.ZN (n_0_0_39), .A1 (n_0_0_94), .A2 (n_0_0_52), .B1 (n_0_0_316), .B2 (n_0_0_127));
OAI22_X1 i_0_0_187 (.ZN (n_0_105), .A1 (sps__n11), .A2 (n_0_0_42), .B1 (n_0_0_356), .B2 (n_0_0_39));
AOI22_X1 i_0_0_186 (.ZN (n_0_0_38), .A1 (n_0_0_358), .A2 (n_0_0_150), .B1 (\n[2] ), .B2 (n_0_0_90));
AOI22_X1 i_0_0_185 (.ZN (n_0_0_37), .A1 (n_0_0_52), .A2 (n_0_0_38), .B1 (n_0_0_316), .B2 (n_0_0_46));
OAI22_X1 i_0_0_184 (.ZN (n_0_104), .A1 (sps__n11), .A2 (n_0_0_41), .B1 (n_0_0_356), .B2 (n_0_0_37));
NOR2_X1 i_0_0_183 (.ZN (n_0_0_36), .A1 (sps__n1), .A2 (n_0_0_340));
AOI22_X1 i_0_0_182 (.ZN (n_0_0_35), .A1 (n_0_0_316), .A2 (n_0_0_110), .B1 (n_0_0_143), .B2 (n_0_0_36));
OAI22_X1 i_0_0_181 (.ZN (n_0_103), .A1 (sps__n11), .A2 (n_0_0_39), .B1 (n_0_0_356), .B2 (n_0_0_35));
AOI22_X1 i_0_0_180 (.ZN (n_0_0_34), .A1 (n_0_0_316), .A2 (n_0_0_101), .B1 (n_0_0_136), .B2 (n_0_0_36));
OAI22_X1 i_0_0_179 (.ZN (n_0_102), .A1 (sps__n11), .A2 (n_0_0_37), .B1 (n_0_0_356), .B2 (n_0_0_34));
AOI22_X1 i_0_0_178 (.ZN (n_0_0_33), .A1 (n_0_0_316), .A2 (n_0_0_94), .B1 (n_0_0_129), .B2 (n_0_0_36));
OAI22_X1 i_0_0_177 (.ZN (n_0_101), .A1 (sps__n11), .A2 (n_0_0_35), .B1 (n_0_0_356), .B2 (n_0_0_33));
AOI22_X1 i_0_0_176 (.ZN (n_0_0_32), .A1 (n_0_0_316), .A2 (n_0_0_38), .B1 (n_0_0_120), .B2 (n_0_0_36));
OAI22_X1 i_0_0_175 (.ZN (n_0_100), .A1 (sps__n11), .A2 (n_0_0_34), .B1 (n_0_0_356), .B2 (n_0_0_32));
AOI22_X1 i_0_0_174 (.ZN (n_0_0_31), .A1 (n_0_0_314), .A2 (n_0_0_143), .B1 (n_0_0_112), .B2 (n_0_0_36));
OAI22_X1 i_0_0_173 (.ZN (n_0_99), .A1 (sps__n11), .A2 (n_0_0_33), .B1 (n_0_0_356), .B2 (n_0_0_31));
AOI22_X1 i_0_0_172 (.ZN (n_0_0_30), .A1 (n_0_0_314), .A2 (n_0_0_136), .B1 (n_0_0_103), .B2 (n_0_0_36));
OAI22_X1 i_0_0_171 (.ZN (n_0_98), .A1 (sps__n11), .A2 (n_0_0_32), .B1 (n_0_0_356), .B2 (n_0_0_30));
AOI22_X1 i_0_0_170 (.ZN (n_0_0_29), .A1 (n_0_0_314), .A2 (n_0_0_129), .B1 (n_0_0_96), .B2 (n_0_0_36));
OAI22_X1 i_0_0_169 (.ZN (n_0_97), .A1 (sps__n11), .A2 (n_0_0_31), .B1 (n_0_0_356), .B2 (n_0_0_29));
NAND2_X1 i_0_0_168 (.ZN (n_0_0_28), .A1 (n_0_0_89), .A2 (n_0_0_36));
OAI21_X1 i_0_0_167 (.ZN (n_0_0_27), .A (n_0_0_28), .B1 (n_0_0_315), .B2 (n_0_0_119));
NAND2_X1 i_0_0_166 (.ZN (n_0_0_26), .A1 (sps__n11), .A2 (n_0_0_27));
OAI21_X1 i_0_0_165 (.ZN (n_0_96), .A (n_0_0_26), .B1 (sps__n11), .B2 (n_0_0_30));
NAND2_X1 i_0_0_164 (.ZN (n_0_0_25), .A1 (n_0_0_338), .A2 (n_0_0_112));
OAI21_X1 i_0_0_163 (.ZN (n_0_95), .A (n_0_0_25), .B1 (sps__n11), .B2 (n_0_0_29));
AOI22_X1 i_0_0_162 (.ZN (n_0_0_24), .A1 (n_0_0_338), .A2 (n_0_0_103), .B1 (n_0_0_356), .B2 (n_0_0_27));
INV_X1 i_0_0_161 (.ZN (n_0_94), .A (n_0_0_24));
NOR2_X1 i_0_0_160 (.ZN (n_0_0_23), .A1 (sps__n11), .A2 (n_0_0_315));
AOI22_X1 i_0_0_159 (.ZN (n_0_0_22), .A1 (n_0_0_338), .A2 (n_0_0_96), .B1 (n_0_0_112), .B2 (n_0_0_23));
INV_X1 i_0_0_158 (.ZN (n_0_93), .A (n_0_0_22));
AOI22_X1 i_0_0_157 (.ZN (n_0_0_21), .A1 (n_0_0_103), .A2 (n_0_0_23), .B1 (n_0_0_338), .B2 (n_0_0_89));
INV_X1 i_0_0_156 (.ZN (n_0_92), .A (n_0_0_21));
AND2_X1 i_0_0_155 (.ZN (n_0_91), .A1 (n_0_0_96), .A2 (n_0_0_23));
AND2_X1 i_0_0_154 (.ZN (n_0_90), .A1 (n_0_0_89), .A2 (n_0_0_23));
OR3_X1 i_0_0_153 (.ZN (n_0_86), .A1 (\n[5] ), .A2 (\n[4] ), .A3 (rst));
NOR2_X1 i_0_0_152 (.ZN (n_0_80), .A1 (rst), .A2 (n_0_0_352));
AOI221_X1 i_0_0_151 (.ZN (n_0_0_20), .A (n_0_0_353), .B1 (sps__n11), .B2 (op2[27])
    , .C1 (n_0_0_356), .C2 (op2[29]));
AOI221_X1 i_0_0_150 (.ZN (n_0_0_19), .A (n_0_0_4), .B1 (n_0_0_356), .B2 (op2[25])
    , .C1 (sps__n10), .C2 (op2[23]));
AOI221_X1 i_0_0_149 (.ZN (n_0_0_18), .A (sps__n10), .B1 (op2[9]), .B2 (n_0_0_353)
    , .C1 (op2[13]), .C2 (n_0_0_4));
AOI221_X1 i_0_0_148 (.ZN (n_0_0_17), .A (n_0_0_356), .B1 (op2[7]), .B2 (n_0_0_353)
    , .C1 (op2[11]), .C2 (n_0_0_4));
OAI33_X1 i_0_0_147 (.ZN (n_0_0_16), .A1 (n_0_0_351), .A2 (n_0_0_19), .A3 (n_0_0_20)
    , .B1 (n_0_0_18), .B2 (n_0_0_17), .B3 (n_0_0_6));
NAND2_X1 i_0_0_146 (.ZN (n_0_0_15), .A1 (n_0_80), .A2 (n_0_0_16));
AOI221_X1 i_0_0_145 (.ZN (n_0_0_14), .A (n_0_0_353), .B1 (n_0_0_356), .B2 (op2[21])
    , .C1 (sps__n11), .C2 (op2[19]));
AOI221_X1 i_0_0_144 (.ZN (n_0_0_13), .A (n_0_0_4), .B1 (n_0_0_356), .B2 (op2[17])
    , .C1 (sps__n11), .C2 (op2[15]));
AOI221_X1 i_0_0_143 (.ZN (n_0_0_12), .A (sps__n10), .B1 (op2[5]), .B2 (n_0_0_4), .C1 (op2[1]), .C2 (n_0_0_353));
AOI221_X1 i_0_0_142 (.ZN (n_0_0_11), .A (n_0_0_356), .B1 (op2[3]), .B2 (n_0_0_4), .C1 (op2[31]), .C2 (n_0_0_353));
OAI33_X1 i_0_0_141 (.ZN (n_0_0_10), .A1 (n_0_0_351), .A2 (n_0_0_13), .A3 (n_0_0_14)
    , .B1 (n_0_0_12), .B2 (n_0_0_11), .B3 (n_0_0_6));
NAND3_X1 i_0_0_140 (.ZN (n_0_0_9), .A1 (n_0_0_354), .A2 (n_0_0_352), .A3 (n_0_0_10));
NAND2_X1 i_0_0_139 (.ZN (n_0_85), .A1 (n_0_0_15), .A2 (n_0_0_9));
OAI21_X1 i_0_0_138 (.ZN (n_0_84), .A (n_0_0_354), .B1 (\n[5] ), .B2 (\n[4] ));
NOR2_X1 i_0_0_137 (.ZN (n_0_0_8), .A1 (\n[5] ), .A2 (n_0_0_3));
AOI211_X1 i_0_0_136 (.ZN (n_0_83), .A (rst), .B (n_0_0_8), .C1 (\n[5] ), .C2 (n_0_0_3));
AND2_X1 i_0_0_135 (.ZN (n_0_82), .A1 (n_0_0_354), .A2 (n_0_0_7));
NOR2_X1 i_0_0_134 (.ZN (n_0_81), .A1 (rst), .A2 (n_0_0_351));
NOR2_X1 i_0_0_133 (.ZN (n_0_79), .A1 (rst), .A2 (n_0_0_353));
NOR2_X1 i_0_0_132 (.ZN (n_0_78), .A1 (sps__n10), .A2 (rst));
AND2_X1 i_0_0_131 (.ZN (n_0_278), .A1 (n_0_0_354), .A2 (n_0_214));
AND2_X1 i_0_0_130 (.ZN (n_0_277), .A1 (n_0_0_354), .A2 (n_0_213));
AND2_X1 i_0_0_129 (.ZN (n_0_276), .A1 (n_0_0_354), .A2 (n_0_212));
AND2_X1 i_0_0_128 (.ZN (n_0_275), .A1 (n_0_0_354), .A2 (n_0_211));
AND2_X1 i_0_0_127 (.ZN (n_0_274), .A1 (n_0_0_354), .A2 (n_0_210));
AND2_X1 i_0_0_126 (.ZN (n_0_273), .A1 (n_0_0_354), .A2 (n_0_209));
AND2_X1 i_0_0_125 (.ZN (n_0_272), .A1 (n_0_0_354), .A2 (n_0_208));
AND2_X1 i_0_0_124 (.ZN (n_0_271), .A1 (n_0_0_354), .A2 (n_0_207));
AND2_X1 i_0_0_123 (.ZN (n_0_270), .A1 (n_0_0_354), .A2 (n_0_206));
AND2_X1 i_0_0_122 (.ZN (n_0_269), .A1 (n_0_0_354), .A2 (n_0_205));
AND2_X1 i_0_0_121 (.ZN (n_0_268), .A1 (n_0_0_354), .A2 (n_0_204));
AND2_X1 i_0_0_120 (.ZN (n_0_267), .A1 (n_0_0_354), .A2 (n_0_203));
AND2_X1 i_0_0_119 (.ZN (n_0_266), .A1 (n_0_0_354), .A2 (n_0_202));
AND2_X1 i_0_0_118 (.ZN (n_0_265), .A1 (n_0_0_354), .A2 (n_0_201));
AND2_X1 i_0_0_117 (.ZN (n_0_264), .A1 (n_0_0_354), .A2 (n_0_200));
AND2_X1 i_0_0_116 (.ZN (n_0_263), .A1 (n_0_0_354), .A2 (n_0_199));
AND2_X1 i_0_0_115 (.ZN (n_0_262), .A1 (n_0_0_354), .A2 (n_0_198));
AND2_X1 i_0_0_114 (.ZN (n_0_261), .A1 (n_0_0_354), .A2 (n_0_197));
AND2_X1 i_0_0_113 (.ZN (n_0_260), .A1 (n_0_0_354), .A2 (n_0_196));
AND2_X1 i_0_0_112 (.ZN (n_0_259), .A1 (n_0_0_354), .A2 (n_0_195));
AND2_X1 i_0_0_111 (.ZN (n_0_258), .A1 (n_0_0_354), .A2 (n_0_194));
AND2_X1 i_0_0_110 (.ZN (n_0_257), .A1 (n_0_0_354), .A2 (n_0_193));
AND2_X1 i_0_0_109 (.ZN (n_0_256), .A1 (n_0_0_354), .A2 (n_0_192));
AND2_X1 i_0_0_108 (.ZN (n_0_255), .A1 (n_0_0_354), .A2 (n_0_191));
AND2_X1 i_0_0_107 (.ZN (n_0_254), .A1 (n_0_0_354), .A2 (n_0_190));
AND2_X1 i_0_0_106 (.ZN (n_0_253), .A1 (n_0_0_354), .A2 (n_0_189));
AND2_X1 i_0_0_105 (.ZN (n_0_252), .A1 (n_0_0_354), .A2 (n_0_188));
AND2_X1 i_0_0_104 (.ZN (n_0_251), .A1 (n_0_0_354), .A2 (n_0_187));
AND2_X1 i_0_0_103 (.ZN (n_0_250), .A1 (n_0_0_354), .A2 (n_0_186));
AND2_X1 i_0_0_102 (.ZN (n_0_249), .A1 (n_0_0_354), .A2 (n_0_185));
AND2_X1 i_0_0_101 (.ZN (n_0_248), .A1 (n_0_0_354), .A2 (n_0_184));
AND2_X1 i_0_0_100 (.ZN (n_0_247), .A1 (n_0_0_354), .A2 (n_0_183));
AND2_X1 i_0_0_99 (.ZN (n_0_246), .A1 (n_0_0_354), .A2 (n_0_182));
AND2_X1 i_0_0_98 (.ZN (n_0_245), .A1 (n_0_0_354), .A2 (n_0_181));
AND2_X1 i_0_0_97 (.ZN (n_0_244), .A1 (n_0_0_354), .A2 (n_0_180));
AND2_X1 i_0_0_96 (.ZN (n_0_243), .A1 (n_0_0_354), .A2 (n_0_179));
AND2_X1 i_0_0_95 (.ZN (n_0_242), .A1 (n_0_0_354), .A2 (n_0_178));
AND2_X1 i_0_0_94 (.ZN (n_0_241), .A1 (n_0_0_354), .A2 (n_0_177));
AND2_X1 i_0_0_93 (.ZN (n_0_240), .A1 (n_0_0_354), .A2 (n_0_176));
AND2_X1 i_0_0_92 (.ZN (n_0_239), .A1 (n_0_0_354), .A2 (n_0_175));
AND2_X1 i_0_0_91 (.ZN (n_0_238), .A1 (n_0_0_354), .A2 (n_0_174));
AND2_X1 i_0_0_90 (.ZN (n_0_237), .A1 (n_0_0_354), .A2 (n_0_173));
AND2_X1 i_0_0_89 (.ZN (n_0_236), .A1 (n_0_0_354), .A2 (n_0_172));
AND2_X1 i_0_0_88 (.ZN (n_0_235), .A1 (n_0_0_354), .A2 (n_0_171));
AND2_X1 i_0_0_87 (.ZN (n_0_234), .A1 (n_0_0_354), .A2 (n_0_170));
AND2_X1 i_0_0_86 (.ZN (n_0_233), .A1 (n_0_0_354), .A2 (n_0_169));
AND2_X1 i_0_0_85 (.ZN (n_0_232), .A1 (n_0_0_354), .A2 (n_0_168));
AND2_X1 i_0_0_84 (.ZN (n_0_231), .A1 (n_0_0_354), .A2 (n_0_167));
AND2_X1 i_0_0_83 (.ZN (n_0_230), .A1 (n_0_0_354), .A2 (n_0_166));
AND2_X1 i_0_0_82 (.ZN (n_0_229), .A1 (n_0_0_354), .A2 (n_0_165));
AND2_X1 i_0_0_81 (.ZN (n_0_228), .A1 (n_0_0_354), .A2 (n_0_164));
AND2_X1 i_0_0_80 (.ZN (n_0_227), .A1 (n_0_0_354), .A2 (n_0_163));
AND2_X1 i_0_0_79 (.ZN (n_0_226), .A1 (n_0_0_354), .A2 (n_0_162));
AND2_X1 i_0_0_78 (.ZN (n_0_225), .A1 (n_0_0_354), .A2 (n_0_161));
AND2_X1 i_0_0_77 (.ZN (n_0_224), .A1 (n_0_0_354), .A2 (n_0_160));
AND2_X1 i_0_0_76 (.ZN (n_0_223), .A1 (n_0_0_354), .A2 (n_0_159));
AND2_X1 i_0_0_75 (.ZN (n_0_222), .A1 (n_0_0_354), .A2 (n_0_158));
AND2_X1 i_0_0_74 (.ZN (n_0_221), .A1 (n_0_0_354), .A2 (n_0_157));
AND2_X1 i_0_0_73 (.ZN (n_0_220), .A1 (n_0_0_354), .A2 (n_0_156));
AND2_X1 i_0_0_72 (.ZN (n_0_219), .A1 (n_0_0_354), .A2 (n_0_155));
AND2_X1 i_0_0_71 (.ZN (n_0_218), .A1 (n_0_0_354), .A2 (n_0_154));
AND2_X1 i_0_0_70 (.ZN (n_0_217), .A1 (n_0_0_354), .A2 (n_0_153));
AND2_X1 i_0_0_69 (.ZN (n_0_216), .A1 (n_0_0_354), .A2 (n_0_152));
AND2_X1 i_0_0_68 (.ZN (n_0_215), .A1 (n_0_0_354), .A2 (n_0_151));
AND2_X1 i_0_0_67 (.ZN (n_0_77), .A1 (n_0_0_354), .A2 (\adder[63] ));
AND2_X1 i_0_0_66 (.ZN (n_0_76), .A1 (n_0_0_354), .A2 (\adder[62] ));
AND2_X1 i_0_0_65 (.ZN (n_0_75), .A1 (n_0_0_354), .A2 (\adder[61] ));
AND2_X1 i_0_0_64 (.ZN (n_0_74), .A1 (n_0_0_354), .A2 (\adder[60] ));
AND2_X1 i_0_0_63 (.ZN (n_0_73), .A1 (n_0_0_354), .A2 (\adder[59] ));
AND2_X1 i_0_0_62 (.ZN (n_0_72), .A1 (n_0_0_354), .A2 (\adder[58] ));
AND2_X1 i_0_0_61 (.ZN (n_0_71), .A1 (n_0_0_354), .A2 (\adder[57] ));
AND2_X1 i_0_0_60 (.ZN (n_0_70), .A1 (n_0_0_354), .A2 (\adder[56] ));
AND2_X1 i_0_0_59 (.ZN (n_0_69), .A1 (n_0_0_354), .A2 (\adder[55] ));
AND2_X1 i_0_0_58 (.ZN (n_0_68), .A1 (n_0_0_354), .A2 (\adder[54] ));
AND2_X1 i_0_0_57 (.ZN (n_0_67), .A1 (n_0_0_354), .A2 (\adder[53] ));
AND2_X1 i_0_0_56 (.ZN (n_0_66), .A1 (n_0_0_354), .A2 (\adder[52] ));
AND2_X1 i_0_0_55 (.ZN (n_0_65), .A1 (n_0_0_354), .A2 (\adder[51] ));
AND2_X1 i_0_0_54 (.ZN (n_0_64), .A1 (n_0_0_354), .A2 (\adder[50] ));
AND2_X1 i_0_0_53 (.ZN (n_0_63), .A1 (n_0_0_354), .A2 (\adder[49] ));
AND2_X1 i_0_0_52 (.ZN (n_0_62), .A1 (n_0_0_354), .A2 (\adder[48] ));
AND2_X1 i_0_0_51 (.ZN (n_0_61), .A1 (n_0_0_354), .A2 (\adder[47] ));
AND2_X1 i_0_0_50 (.ZN (n_0_60), .A1 (n_0_0_354), .A2 (\adder[46] ));
AND2_X1 i_0_0_49 (.ZN (n_0_59), .A1 (n_0_0_354), .A2 (\adder[45] ));
AND2_X1 i_0_0_48 (.ZN (n_0_58), .A1 (n_0_0_354), .A2 (\adder[44] ));
AND2_X1 i_0_0_47 (.ZN (n_0_57), .A1 (n_0_0_354), .A2 (\adder[43] ));
AND2_X1 i_0_0_46 (.ZN (n_0_56), .A1 (n_0_0_354), .A2 (\adder[42] ));
AND2_X1 i_0_0_45 (.ZN (n_0_55), .A1 (n_0_0_354), .A2 (\adder[41] ));
AND2_X1 i_0_0_44 (.ZN (n_0_54), .A1 (n_0_0_354), .A2 (\adder[40] ));
AND2_X1 i_0_0_43 (.ZN (n_0_53), .A1 (n_0_0_354), .A2 (\adder[39] ));
AND2_X1 i_0_0_42 (.ZN (n_0_52), .A1 (n_0_0_354), .A2 (\adder[38] ));
AND2_X1 i_0_0_41 (.ZN (n_0_51), .A1 (n_0_0_354), .A2 (\adder[37] ));
AND2_X1 i_0_0_40 (.ZN (n_0_50), .A1 (n_0_0_354), .A2 (\adder[36] ));
AND2_X1 i_0_0_39 (.ZN (n_0_49), .A1 (n_0_0_354), .A2 (\adder[35] ));
AND2_X1 i_0_0_38 (.ZN (n_0_48), .A1 (n_0_0_354), .A2 (\adder[34] ));
AND2_X1 i_0_0_37 (.ZN (n_0_47), .A1 (n_0_0_354), .A2 (\adder[33] ));
AND2_X1 i_0_0_36 (.ZN (n_0_46), .A1 (n_0_0_354), .A2 (\adder[32] ));
AND2_X1 i_0_0_35 (.ZN (n_0_45), .A1 (n_0_0_354), .A2 (\adder[31] ));
AND2_X1 i_0_0_34 (.ZN (n_0_44), .A1 (n_0_0_354), .A2 (\adder[30] ));
AND2_X1 i_0_0_33 (.ZN (n_0_43), .A1 (n_0_0_354), .A2 (\adder[29] ));
AND2_X1 i_0_0_32 (.ZN (n_0_42), .A1 (n_0_0_354), .A2 (\adder[28] ));
AND2_X1 i_0_0_31 (.ZN (n_0_41), .A1 (n_0_0_354), .A2 (\adder[27] ));
AND2_X1 i_0_0_30 (.ZN (n_0_40), .A1 (n_0_0_354), .A2 (\adder[26] ));
AND2_X1 i_0_0_29 (.ZN (n_0_39), .A1 (n_0_0_354), .A2 (\adder[25] ));
AND2_X1 i_0_0_28 (.ZN (n_0_38), .A1 (n_0_0_354), .A2 (\adder[24] ));
AND2_X1 i_0_0_27 (.ZN (n_0_37), .A1 (n_0_0_354), .A2 (\adder[23] ));
AND2_X1 i_0_0_26 (.ZN (n_0_36), .A1 (n_0_0_354), .A2 (\adder[22] ));
AND2_X1 i_0_0_25 (.ZN (n_0_35), .A1 (n_0_0_354), .A2 (\adder[21] ));
AND2_X1 i_0_0_24 (.ZN (n_0_34), .A1 (n_0_0_354), .A2 (\adder[20] ));
AND2_X1 i_0_0_23 (.ZN (n_0_2), .A1 (n_0_0_354), .A2 (\adder[19] ));
AND2_X1 i_0_0_22 (.ZN (n_0_1), .A1 (n_0_0_354), .A2 (\adder[18] ));
AND2_X1 i_0_0_21 (.ZN (n_0_296), .A1 (n_0_0_354), .A2 (\adder[17] ));
AND2_X1 i_0_0_20 (.ZN (n_0_295), .A1 (n_0_0_354), .A2 (\adder[16] ));
AND2_X1 i_0_0_19 (.ZN (n_0_294), .A1 (n_0_0_354), .A2 (\adder[15] ));
AND2_X1 i_0_0_18 (.ZN (n_0_293), .A1 (n_0_0_354), .A2 (\adder[14] ));
AND2_X1 i_0_0_17 (.ZN (n_0_292), .A1 (n_0_0_354), .A2 (\adder[13] ));
AND2_X1 i_0_0_16 (.ZN (n_0_291), .A1 (n_0_0_354), .A2 (\adder[12] ));
AND2_X1 i_0_0_15 (.ZN (n_0_290), .A1 (n_0_0_354), .A2 (\adder[11] ));
AND2_X1 i_0_0_14 (.ZN (n_0_289), .A1 (n_0_0_354), .A2 (\adder[10] ));
AND2_X1 i_0_0_13 (.ZN (n_0_288), .A1 (n_0_0_354), .A2 (\adder[9] ));
AND2_X1 i_0_0_12 (.ZN (n_0_287), .A1 (n_0_0_354), .A2 (\adder[8] ));
AND2_X1 i_0_0_11 (.ZN (n_0_286), .A1 (n_0_0_354), .A2 (\adder[7] ));
AND2_X1 i_0_0_10 (.ZN (n_0_285), .A1 (n_0_0_354), .A2 (\adder[6] ));
AND2_X1 i_0_0_9 (.ZN (n_0_284), .A1 (n_0_0_354), .A2 (\adder[5] ));
AND2_X1 i_0_0_8 (.ZN (n_0_283), .A1 (n_0_0_354), .A2 (\adder[4] ));
AND2_X1 i_0_0_7 (.ZN (n_0_282), .A1 (n_0_0_354), .A2 (\adder[3] ));
AND2_X1 i_0_0_6 (.ZN (n_0_281), .A1 (n_0_0_354), .A2 (\adder[2] ));
AND2_X1 i_0_0_5 (.ZN (n_0_280), .A1 (n_0_0_354), .A2 (\adder[1] ));
AND2_X1 i_0_0_4 (.ZN (n_0_279), .A1 (n_0_0_354), .A2 (\adder[0] ));
HA_X1 i_0_0_3 (.CO (n_0_0_3), .S (n_0_0_7), .A (\n[4] ), .B (n_0_0_2));
HA_X1 i_0_0_2 (.CO (n_0_0_2), .S (n_0_0_6), .A (\n[3] ), .B (n_0_0_1));
HA_X1 i_0_0_1 (.CO (n_0_0_1), .S (n_0_0_5), .A (\n[2] ), .B (n_0_0_0));
HA_X1 i_0_0_0 (.CO (n_0_0_0), .S (n_0_0_4), .A (sps__n7), .B (sps__n11));
datapath__0_16 i_0_14 (.p_1 ({n_0_214, n_0_213, n_0_212, n_0_211, n_0_210, n_0_209, 
    n_0_208, n_0_207, n_0_206, n_0_205, n_0_204, n_0_203, n_0_202, n_0_201, n_0_200, 
    n_0_199, n_0_198, n_0_197, n_0_196, n_0_195, n_0_194, n_0_193, n_0_192, n_0_191, 
    n_0_190, n_0_189, n_0_188, n_0_187, n_0_186, n_0_185, n_0_184, n_0_183, n_0_182, 
    n_0_181, n_0_180, n_0_179, n_0_178, n_0_177, n_0_176, n_0_175, n_0_174, n_0_173, 
    n_0_172, n_0_171, n_0_170, n_0_169, n_0_168, n_0_167, n_0_166, n_0_165, n_0_164, 
    n_0_163, n_0_162, n_0_161, n_0_160, n_0_159, n_0_158, n_0_157, n_0_156, n_0_155, 
    n_0_154, n_0_153, n_0_152, n_0_151}), .adder ({\adder[63] , \adder[62] , \adder[61] , 
    \adder[60] , \adder[59] , \adder[58] , \adder[57] , \adder[56] , \adder[55] , 
    \adder[54] , \adder[53] , \adder[52] , \adder[51] , \adder[50] , \adder[49] , 
    \adder[48] , \adder[47] , \adder[46] , \adder[45] , \adder[44] , \adder[43] , 
    \adder[42] , \adder[41] , \adder[40] , \adder[39] , \adder[38] , \adder[37] , 
    \adder[36] , \adder[35] , \adder[34] , \adder[33] , \adder[32] , \adder[31] , 
    \adder[30] , \adder[29] , \adder[28] , \adder[27] , \adder[26] , \adder[25] , 
    \adder[24] , \adder[23] , \adder[22] , \adder[21] , \adder[20] , \adder[19] , 
    \adder[18] , \adder[17] , \adder[16] , \adder[15] , \adder[14] , \adder[13] , 
    \adder[12] , \adder[11] , \adder[10] , \adder[9] , \adder[8] , \adder[7] , \adder[6] , 
    \adder[5] , \adder[4] , \adder[3] , \adder[2] , \adder[1] , \adder[0] }), .p_0 ({
    uc_1, uc_2, n_0_89, n_0_150, n_0_149, n_0_148, n_0_147, n_0_146, n_0_145, n_0_144, 
    n_0_143, n_0_142, n_0_141, n_0_140, n_0_139, n_0_138, n_0_137, n_0_136, n_0_135, 
    n_0_134, n_0_133, n_0_132, n_0_131, n_0_130, n_0_129, n_0_128, n_0_127, n_0_126, 
    n_0_125, n_0_124, n_0_123, n_0_122, n_0_121, n_0_120, n_0_119, n_0_118, n_0_117, 
    n_0_116, n_0_115, n_0_114, n_0_113, n_0_112, n_0_111, n_0_110, n_0_109, n_0_108, 
    n_0_107, n_0_106, n_0_105, n_0_104, n_0_103, n_0_102, n_0_101, n_0_100, n_0_99, 
    n_0_98, n_0_97, n_0_96, n_0_95, n_0_94, n_0_93, n_0_92, n_0_91, n_0_90}));
datapath i_0_2 (.p_0 ({n_0_33, n_0_32, n_0_31, n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, 
    n_0_25, n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, 
    n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, n_0_5, 
    n_0_4, n_0_3, uc_0}), .op1 ({op1[31], op1[30], op1[29], op1[28], op1[27], op1[26], 
    op1[25], op1[24], op1[23], op1[22], op1[21], op1[20], op1[19], op1[18], op1[17], 
    op1[16], op1[15], op1[14], op1[13], op1[12], op1[11], op1[10], op1[9], op1[8], 
    op1[7], op1[6], op1[5], op1[4], op1[3], op1[2], op1[1], op1[0]}));
DFF_X1 \P_reg[0]  (.Q (P[0]), .CK (n_0_0), .D (n_0_279));
DFF_X1 \P_reg[1]  (.Q (P[1]), .CK (n_0_0), .D (n_0_280));
DFF_X1 \P_reg[2]  (.Q (P[2]), .CK (n_0_0), .D (n_0_281));
DFF_X1 \P_reg[3]  (.Q (P[3]), .CK (n_0_0), .D (n_0_282));
DFF_X1 \P_reg[4]  (.Q (P[4]), .CK (n_0_0), .D (n_0_283));
DFF_X1 \P_reg[5]  (.Q (P[5]), .CK (n_0_0), .D (n_0_284));
DFF_X1 \P_reg[6]  (.Q (P[6]), .CK (n_0_0), .D (n_0_285));
DFF_X1 \P_reg[7]  (.Q (P[7]), .CK (n_0_0), .D (n_0_286));
DFF_X1 \P_reg[8]  (.Q (P[8]), .CK (n_0_0), .D (n_0_287));
DFF_X1 \P_reg[9]  (.Q (P[9]), .CK (n_0_0), .D (n_0_288));
DFF_X1 \P_reg[10]  (.Q (P[10]), .CK (n_0_0), .D (n_0_289));
DFF_X1 \P_reg[11]  (.Q (P[11]), .CK (n_0_0), .D (n_0_290));
DFF_X1 \P_reg[12]  (.Q (P[12]), .CK (n_0_0), .D (n_0_291));
DFF_X1 \P_reg[13]  (.Q (P[13]), .CK (n_0_0), .D (n_0_292));
DFF_X1 \P_reg[14]  (.Q (P[14]), .CK (n_0_0), .D (n_0_293));
DFF_X1 \P_reg[15]  (.Q (P[15]), .CK (n_0_0), .D (n_0_294));
DFF_X1 \P_reg[16]  (.Q (P[16]), .CK (n_0_0), .D (n_0_295));
DFF_X1 \P_reg[17]  (.Q (P[17]), .CK (n_0_0), .D (n_0_296));
DFF_X1 \P_reg[18]  (.Q (P[18]), .CK (n_0_0), .D (n_0_1));
DFF_X1 \P_reg[19]  (.Q (P[19]), .CK (n_0_0), .D (n_0_2));
DFF_X1 \P_reg[20]  (.Q (P[20]), .CK (n_0_0), .D (n_0_34));
DFF_X1 \P_reg[21]  (.Q (P[21]), .CK (n_0_0), .D (n_0_35));
DFF_X1 \P_reg[22]  (.Q (P[22]), .CK (n_0_0), .D (n_0_36));
DFF_X1 \P_reg[23]  (.Q (P[23]), .CK (n_0_0), .D (n_0_37));
DFF_X1 \P_reg[24]  (.Q (P[24]), .CK (n_0_0), .D (n_0_38));
DFF_X1 \P_reg[25]  (.Q (P[25]), .CK (n_0_0), .D (n_0_39));
DFF_X1 \P_reg[26]  (.Q (P[26]), .CK (n_0_0), .D (n_0_40));
DFF_X1 \P_reg[27]  (.Q (P[27]), .CK (n_0_0), .D (n_0_41));
DFF_X1 \P_reg[28]  (.Q (P[28]), .CK (n_0_0), .D (n_0_42));
DFF_X1 \P_reg[29]  (.Q (P[29]), .CK (n_0_0), .D (n_0_43));
DFF_X1 \P_reg[30]  (.Q (P[30]), .CK (n_0_0), .D (n_0_44));
DFF_X1 \P_reg[31]  (.Q (P[31]), .CK (n_0_0), .D (n_0_45));
DFF_X1 \P_reg[32]  (.Q (P[32]), .CK (n_0_0), .D (n_0_46));
DFF_X1 \P_reg[33]  (.Q (P[33]), .CK (n_0_0), .D (n_0_47));
DFF_X1 \P_reg[34]  (.Q (P[34]), .CK (n_0_0), .D (n_0_48));
DFF_X1 \P_reg[35]  (.Q (P[35]), .CK (n_0_0), .D (n_0_49));
DFF_X1 \P_reg[36]  (.Q (P[36]), .CK (n_0_0), .D (n_0_50));
DFF_X1 \P_reg[37]  (.Q (P[37]), .CK (n_0_0), .D (n_0_51));
DFF_X1 \P_reg[38]  (.Q (P[38]), .CK (n_0_0), .D (n_0_52));
DFF_X1 \P_reg[39]  (.Q (P[39]), .CK (n_0_0), .D (n_0_53));
DFF_X1 \P_reg[40]  (.Q (P[40]), .CK (n_0_0), .D (n_0_54));
DFF_X1 \P_reg[41]  (.Q (P[41]), .CK (n_0_0), .D (n_0_55));
DFF_X1 \P_reg[42]  (.Q (P[42]), .CK (n_0_0), .D (n_0_56));
DFF_X1 \P_reg[43]  (.Q (P[43]), .CK (n_0_0), .D (n_0_57));
DFF_X1 \P_reg[44]  (.Q (P[44]), .CK (n_0_0), .D (n_0_58));
DFF_X1 \P_reg[45]  (.Q (P[45]), .CK (n_0_0), .D (n_0_59));
DFF_X1 \P_reg[46]  (.Q (P[46]), .CK (n_0_0), .D (n_0_60));
DFF_X1 \P_reg[47]  (.Q (P[47]), .CK (n_0_0), .D (n_0_61));
DFF_X1 \P_reg[48]  (.Q (P[48]), .CK (n_0_0), .D (n_0_62));
DFF_X1 \P_reg[49]  (.Q (P[49]), .CK (n_0_0), .D (n_0_63));
DFF_X1 \P_reg[50]  (.Q (P[50]), .CK (n_0_0), .D (n_0_64));
DFF_X1 \P_reg[51]  (.Q (P[51]), .CK (n_0_0), .D (n_0_65));
DFF_X1 \P_reg[52]  (.Q (P[52]), .CK (n_0_0), .D (n_0_66));
DFF_X1 \P_reg[53]  (.Q (P[53]), .CK (n_0_0), .D (n_0_67));
DFF_X1 \P_reg[54]  (.Q (P[54]), .CK (n_0_0), .D (n_0_68));
DFF_X1 \P_reg[55]  (.Q (P[55]), .CK (n_0_0), .D (n_0_69));
DFF_X1 \P_reg[56]  (.Q (P[56]), .CK (n_0_0), .D (n_0_70));
DFF_X1 \P_reg[57]  (.Q (P[57]), .CK (n_0_0), .D (n_0_71));
DFF_X1 \P_reg[58]  (.Q (P[58]), .CK (n_0_0), .D (n_0_72));
DFF_X1 \P_reg[59]  (.Q (P[59]), .CK (n_0_0), .D (n_0_73));
DFF_X1 \P_reg[60]  (.Q (P[60]), .CK (n_0_0), .D (n_0_74));
DFF_X1 \P_reg[61]  (.Q (P[61]), .CK (n_0_0), .D (n_0_75));
DFF_X1 \P_reg[62]  (.Q (P[62]), .CK (n_0_0), .D (n_0_76));
DFF_X1 \P_reg[63]  (.Q (P[63]), .CK (n_0_0), .D (n_0_77));
CLKGATETST_X1 clk_gate_P_reg (.GCK (n_0_0), .CK (clk), .E (n_0_86), .SE (1'b0 ));
BUF_X8 sps__L1_c1 (.Z (sps__n1), .A (n_0_0_357));
BUF_X4 sps__L1_c4 (.Z (sps__n4), .A (n_0_0_303));
BUF_X8 sps__L1_c7 (.Z (sps__n7), .A (\n[1] ));
CLKBUF_X3 sps__L1_c10 (.Z (sps__n10), .A (\n[0] ));
BUF_X8 sps__L1_c11 (.Z (sps__n11), .A (\n[0] ));
BUF_X4 sps__L1_c16 (.Z (sps__n16), .A (n_0_0_302));
BUF_X8 spc__L1_c19 (.Z (spc__n19), .A (n_0_0_304));
BUF_X8 spc__L1_c22 (.Z (spc__n22), .A (n_0_0_305));
BUF_X4 spt__c25 (.Z (\n[2] ), .A (spt__n25));

endmodule //Radix4_Booth_new


