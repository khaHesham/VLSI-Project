/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Fri Dec 23 14:56:16 2022
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 1769545571 */

module datapath(A, p_0, M);
   input [31:0]A;
   output [31:0]p_0;
   input [31:0]M;

   INV_X1 i_0 (.A(A[0]), .ZN(n_0));
   NAND2_X1 i_1 (.A1(n_0), .A2(M[0]), .ZN(n_1));
   OAI21_X1 i_2 (.A(n_1), .B1(M[0]), .B2(n_0), .ZN(p_0[0]));
   XNOR2_X1 i_3 (.A(A[1]), .B(M[1]), .ZN(n_2));
   XOR2_X1 i_4 (.A(n_2), .B(n_1), .Z(p_0[1]));
   INV_X1 i_5 (.A(n_1), .ZN(n_3));
   INV_X1 i_6 (.A(A[1]), .ZN(n_4));
   AOI22_X1 i_7 (.A1(n_2), .A2(n_3), .B1(n_4), .B2(M[1]), .ZN(n_5));
   XOR2_X1 i_8 (.A(M[2]), .B(A[2]), .Z(n_6));
   XNOR2_X1 i_9 (.A(n_5), .B(n_6), .ZN(p_0[2]));
   INV_X1 i_10 (.A(M[2]), .ZN(n_7));
   OAI22_X1 i_11 (.A1(n_5), .A2(n_6), .B1(n_7), .B2(A[2]), .ZN(n_8));
   XNOR2_X1 i_12 (.A(A[3]), .B(M[3]), .ZN(n_9));
   XNOR2_X1 i_13 (.A(n_8), .B(n_9), .ZN(p_0[3]));
   INV_X1 i_14 (.A(A[3]), .ZN(n_10));
   AOI22_X1 i_15 (.A1(n_8), .A2(n_9), .B1(n_10), .B2(M[3]), .ZN(n_11));
   XOR2_X1 i_16 (.A(A[4]), .B(M[4]), .Z(n_12));
   XNOR2_X1 i_17 (.A(n_11), .B(n_12), .ZN(p_0[4]));
   INV_X1 i_18 (.A(M[4]), .ZN(n_13));
   OAI22_X1 i_19 (.A1(n_11), .A2(n_12), .B1(n_13), .B2(A[4]), .ZN(n_14));
   XNOR2_X1 i_20 (.A(A[5]), .B(M[5]), .ZN(n_15));
   XNOR2_X1 i_21 (.A(n_14), .B(n_15), .ZN(p_0[5]));
   INV_X1 i_22 (.A(A[5]), .ZN(n_16));
   AOI22_X1 i_23 (.A1(n_14), .A2(n_15), .B1(n_16), .B2(M[5]), .ZN(n_17));
   XOR2_X1 i_24 (.A(A[6]), .B(M[6]), .Z(n_18));
   XNOR2_X1 i_25 (.A(n_17), .B(n_18), .ZN(p_0[6]));
   INV_X1 i_26 (.A(M[6]), .ZN(n_19));
   OAI22_X1 i_27 (.A1(n_17), .A2(n_18), .B1(n_19), .B2(A[6]), .ZN(n_20));
   XNOR2_X1 i_28 (.A(A[7]), .B(M[7]), .ZN(n_21));
   XNOR2_X1 i_29 (.A(n_20), .B(n_21), .ZN(p_0[7]));
   INV_X1 i_30 (.A(A[7]), .ZN(n_22));
   AOI22_X1 i_31 (.A1(n_20), .A2(n_21), .B1(n_22), .B2(M[7]), .ZN(n_23));
   XOR2_X1 i_32 (.A(A[8]), .B(M[8]), .Z(n_24));
   XNOR2_X1 i_33 (.A(n_23), .B(n_24), .ZN(p_0[8]));
   INV_X1 i_34 (.A(M[8]), .ZN(n_25));
   OAI22_X1 i_35 (.A1(n_23), .A2(n_24), .B1(n_25), .B2(A[8]), .ZN(n_26));
   XNOR2_X1 i_36 (.A(A[9]), .B(M[9]), .ZN(n_27));
   XNOR2_X1 i_37 (.A(n_26), .B(n_27), .ZN(p_0[9]));
   INV_X1 i_38 (.A(A[9]), .ZN(n_28));
   AOI22_X1 i_39 (.A1(n_26), .A2(n_27), .B1(n_28), .B2(M[9]), .ZN(n_29));
   XOR2_X1 i_40 (.A(A[10]), .B(M[10]), .Z(n_30));
   XNOR2_X1 i_41 (.A(n_29), .B(n_30), .ZN(p_0[10]));
   INV_X1 i_42 (.A(M[10]), .ZN(n_31));
   OAI22_X1 i_43 (.A1(n_29), .A2(n_30), .B1(n_31), .B2(A[10]), .ZN(n_32));
   XNOR2_X1 i_44 (.A(A[11]), .B(M[11]), .ZN(n_33));
   XNOR2_X1 i_45 (.A(n_32), .B(n_33), .ZN(p_0[11]));
   INV_X1 i_46 (.A(A[11]), .ZN(n_34));
   AOI22_X1 i_47 (.A1(n_32), .A2(n_33), .B1(n_34), .B2(M[11]), .ZN(n_35));
   XOR2_X1 i_48 (.A(A[12]), .B(M[12]), .Z(n_36));
   XNOR2_X1 i_49 (.A(n_35), .B(n_36), .ZN(p_0[12]));
   INV_X1 i_50 (.A(M[12]), .ZN(n_37));
   OAI22_X1 i_51 (.A1(n_35), .A2(n_36), .B1(n_37), .B2(A[12]), .ZN(n_38));
   XNOR2_X1 i_52 (.A(A[13]), .B(M[13]), .ZN(n_39));
   XNOR2_X1 i_53 (.A(n_38), .B(n_39), .ZN(p_0[13]));
   INV_X1 i_54 (.A(A[13]), .ZN(n_40));
   AOI22_X1 i_55 (.A1(n_38), .A2(n_39), .B1(n_40), .B2(M[13]), .ZN(n_41));
   XOR2_X1 i_56 (.A(A[14]), .B(M[14]), .Z(n_42));
   XNOR2_X1 i_57 (.A(n_41), .B(n_42), .ZN(p_0[14]));
   INV_X1 i_58 (.A(M[14]), .ZN(n_43));
   OAI22_X1 i_59 (.A1(n_41), .A2(n_42), .B1(n_43), .B2(A[14]), .ZN(n_44));
   XNOR2_X1 i_60 (.A(A[15]), .B(M[15]), .ZN(n_45));
   XNOR2_X1 i_61 (.A(n_44), .B(n_45), .ZN(p_0[15]));
   INV_X1 i_62 (.A(A[15]), .ZN(n_46));
   AOI22_X1 i_63 (.A1(n_44), .A2(n_45), .B1(n_46), .B2(M[15]), .ZN(n_47));
   XOR2_X1 i_64 (.A(A[16]), .B(M[16]), .Z(n_48));
   XNOR2_X1 i_65 (.A(n_47), .B(n_48), .ZN(p_0[16]));
   INV_X1 i_66 (.A(M[16]), .ZN(n_49));
   OAI22_X1 i_67 (.A1(n_47), .A2(n_48), .B1(n_49), .B2(A[16]), .ZN(n_50));
   XNOR2_X1 i_68 (.A(A[17]), .B(M[17]), .ZN(n_51));
   XNOR2_X1 i_69 (.A(n_50), .B(n_51), .ZN(p_0[17]));
   INV_X1 i_70 (.A(A[17]), .ZN(n_52));
   AOI22_X1 i_71 (.A1(n_50), .A2(n_51), .B1(n_52), .B2(M[17]), .ZN(n_53));
   XOR2_X1 i_72 (.A(A[18]), .B(M[18]), .Z(n_54));
   XNOR2_X1 i_73 (.A(n_53), .B(n_54), .ZN(p_0[18]));
   INV_X1 i_74 (.A(M[18]), .ZN(n_55));
   OAI22_X1 i_75 (.A1(n_53), .A2(n_54), .B1(n_55), .B2(A[18]), .ZN(n_56));
   XNOR2_X1 i_76 (.A(A[19]), .B(M[19]), .ZN(n_57));
   XNOR2_X1 i_77 (.A(n_56), .B(n_57), .ZN(p_0[19]));
   INV_X1 i_78 (.A(A[19]), .ZN(n_58));
   AOI22_X1 i_79 (.A1(n_56), .A2(n_57), .B1(n_58), .B2(M[19]), .ZN(n_59));
   XOR2_X1 i_80 (.A(A[20]), .B(M[20]), .Z(n_60));
   XNOR2_X1 i_81 (.A(n_59), .B(n_60), .ZN(p_0[20]));
   INV_X1 i_82 (.A(M[20]), .ZN(n_61));
   OAI22_X1 i_83 (.A1(n_59), .A2(n_60), .B1(n_61), .B2(A[20]), .ZN(n_62));
   XNOR2_X1 i_84 (.A(A[21]), .B(M[21]), .ZN(n_63));
   XNOR2_X1 i_85 (.A(n_62), .B(n_63), .ZN(p_0[21]));
   INV_X1 i_86 (.A(A[21]), .ZN(n_64));
   AOI22_X1 i_87 (.A1(n_62), .A2(n_63), .B1(n_64), .B2(M[21]), .ZN(n_65));
   XOR2_X1 i_88 (.A(A[22]), .B(M[22]), .Z(n_66));
   XNOR2_X1 i_89 (.A(n_65), .B(n_66), .ZN(p_0[22]));
   INV_X1 i_90 (.A(M[22]), .ZN(n_67));
   OAI22_X1 i_91 (.A1(n_65), .A2(n_66), .B1(n_67), .B2(A[22]), .ZN(n_68));
   XNOR2_X1 i_92 (.A(A[23]), .B(M[23]), .ZN(n_69));
   XNOR2_X1 i_93 (.A(n_68), .B(n_69), .ZN(p_0[23]));
   INV_X1 i_94 (.A(A[23]), .ZN(n_70));
   AOI22_X1 i_95 (.A1(n_68), .A2(n_69), .B1(n_70), .B2(M[23]), .ZN(n_71));
   XOR2_X1 i_96 (.A(A[24]), .B(M[24]), .Z(n_72));
   XNOR2_X1 i_97 (.A(n_71), .B(n_72), .ZN(p_0[24]));
   INV_X1 i_98 (.A(M[24]), .ZN(n_73));
   OAI22_X1 i_99 (.A1(n_71), .A2(n_72), .B1(n_73), .B2(A[24]), .ZN(n_74));
   XNOR2_X1 i_100 (.A(A[25]), .B(M[25]), .ZN(n_75));
   XNOR2_X1 i_101 (.A(n_74), .B(n_75), .ZN(p_0[25]));
   INV_X1 i_102 (.A(A[25]), .ZN(n_76));
   AOI22_X1 i_103 (.A1(n_74), .A2(n_75), .B1(n_76), .B2(M[25]), .ZN(n_77));
   XOR2_X1 i_104 (.A(A[26]), .B(M[26]), .Z(n_78));
   XNOR2_X1 i_105 (.A(n_77), .B(n_78), .ZN(p_0[26]));
   INV_X1 i_106 (.A(M[26]), .ZN(n_79));
   OAI22_X1 i_107 (.A1(n_77), .A2(n_78), .B1(n_79), .B2(A[26]), .ZN(n_80));
   XNOR2_X1 i_108 (.A(A[27]), .B(M[27]), .ZN(n_81));
   XNOR2_X1 i_109 (.A(n_80), .B(n_81), .ZN(p_0[27]));
   INV_X1 i_110 (.A(A[27]), .ZN(n_82));
   AOI22_X1 i_111 (.A1(n_80), .A2(n_81), .B1(n_82), .B2(M[27]), .ZN(n_83));
   XOR2_X1 i_112 (.A(A[28]), .B(M[28]), .Z(n_84));
   XNOR2_X1 i_113 (.A(n_83), .B(n_84), .ZN(p_0[28]));
   INV_X1 i_114 (.A(M[28]), .ZN(n_85));
   OAI22_X1 i_115 (.A1(n_83), .A2(n_84), .B1(n_85), .B2(A[28]), .ZN(n_86));
   XNOR2_X1 i_116 (.A(A[29]), .B(M[29]), .ZN(n_87));
   XNOR2_X1 i_117 (.A(n_86), .B(n_87), .ZN(p_0[29]));
   INV_X1 i_118 (.A(A[29]), .ZN(n_88));
   AOI22_X1 i_119 (.A1(n_86), .A2(n_87), .B1(n_88), .B2(M[29]), .ZN(n_89));
   INV_X1 i_120 (.A(A[31]), .ZN(n_90));
   INV_X1 i_121 (.A(M[30]), .ZN(n_91));
   AOI22_X1 i_122 (.A1(n_90), .A2(n_91), .B1(A[31]), .B2(M[30]), .ZN(n_92));
   XNOR2_X1 i_123 (.A(n_89), .B(n_92), .ZN(p_0[30]));
   INV_X1 i_124 (.A(n_89), .ZN(n_93));
   OAI33_X1 i_125 (.A1(n_93), .A2(A[31]), .A3(M[30]), .B1(n_89), .B2(n_90), 
      .B3(n_91), .ZN(n_94));
   XNOR2_X1 i_126 (.A(n_94), .B(M[31]), .ZN(p_0[31]));
endmodule

module datapath__0_1(M, A, p_0);
   input [31:0]M;
   input [31:0]A;
   output [31:0]p_0;

   INV_X1 i_0 (.A(n_0), .ZN(p_0[0]));
   OAI21_X1 i_1 (.A(n_154), .B1(M[0]), .B2(A[0]), .ZN(n_0));
   XOR2_X1 i_2 (.A(n_154), .B(n_1), .Z(p_0[1]));
   OAI21_X1 i_3 (.A(n_153), .B1(M[1]), .B2(A[1]), .ZN(n_1));
   XNOR2_X1 i_4 (.A(n_152), .B(n_2), .ZN(p_0[2]));
   OAI21_X1 i_5 (.A(n_157), .B1(M[2]), .B2(A[2]), .ZN(n_2));
   XOR2_X1 i_6 (.A(n_151), .B(n_3), .Z(p_0[3]));
   OAI21_X1 i_7 (.A(n_158), .B1(n_164), .B2(n_161), .ZN(n_3));
   XOR2_X1 i_8 (.A(n_149), .B(n_10), .Z(p_0[4]));
   XOR2_X1 i_9 (.A(n_9), .B(n_6), .Z(p_0[5]));
   XOR2_X1 i_10 (.A(n_7), .B(n_4), .Z(p_0[6]));
   NOR2_X1 i_11 (.A1(n_146), .A2(n_137), .ZN(n_4));
   XNOR2_X1 i_12 (.A(n_11), .B(n_5), .ZN(p_0[7]));
   OAI22_X1 i_13 (.A1(M[6]), .A2(A[6]), .B1(n_137), .B2(n_7), .ZN(n_5));
   AOI21_X1 i_14 (.A(n_147), .B1(M[5]), .B2(A[5]), .ZN(n_6));
   AOI21_X1 i_15 (.A(n_147), .B1(n_141), .B2(n_8), .ZN(n_7));
   INV_X1 i_16 (.A(n_9), .ZN(n_8));
   AOI21_X1 i_17 (.A(n_144), .B1(n_149), .B2(n_142), .ZN(n_9));
   OAI21_X1 i_18 (.A(n_142), .B1(M[4]), .B2(A[4]), .ZN(n_10));
   NOR2_X1 i_19 (.A1(n_148), .A2(n_139), .ZN(n_11));
   XNOR2_X1 i_20 (.A(n_135), .B(n_18), .ZN(p_0[8]));
   XOR2_X1 i_21 (.A(n_17), .B(n_14), .Z(p_0[9]));
   XOR2_X1 i_22 (.A(n_15), .B(n_12), .Z(p_0[10]));
   NOR2_X1 i_23 (.A1(n_132), .A2(n_123), .ZN(n_12));
   XNOR2_X1 i_24 (.A(n_19), .B(n_13), .ZN(p_0[11]));
   OAI22_X1 i_25 (.A1(M[10]), .A2(A[10]), .B1(n_123), .B2(n_15), .ZN(n_13));
   AOI21_X1 i_26 (.A(n_133), .B1(M[9]), .B2(A[9]), .ZN(n_14));
   AOI21_X1 i_27 (.A(n_133), .B1(n_127), .B2(n_16), .ZN(n_15));
   INV_X1 i_28 (.A(n_17), .ZN(n_16));
   AOI21_X1 i_29 (.A(n_130), .B1(n_135), .B2(n_128), .ZN(n_17));
   AOI21_X1 i_30 (.A(n_130), .B1(M[8]), .B2(A[8]), .ZN(n_18));
   NOR2_X1 i_31 (.A1(n_134), .A2(n_125), .ZN(n_19));
   XOR2_X1 i_32 (.A(n_121), .B(n_26), .Z(p_0[12]));
   XOR2_X1 i_33 (.A(n_25), .B(n_22), .Z(p_0[13]));
   XOR2_X1 i_34 (.A(n_23), .B(n_20), .Z(p_0[14]));
   NOR2_X1 i_35 (.A1(n_118), .A2(n_109), .ZN(n_20));
   XNOR2_X1 i_36 (.A(n_27), .B(n_21), .ZN(p_0[15]));
   OAI22_X1 i_37 (.A1(M[14]), .A2(A[14]), .B1(n_109), .B2(n_23), .ZN(n_21));
   AOI21_X1 i_38 (.A(n_119), .B1(M[13]), .B2(A[13]), .ZN(n_22));
   AOI21_X1 i_39 (.A(n_119), .B1(n_113), .B2(n_24), .ZN(n_23));
   INV_X1 i_40 (.A(n_25), .ZN(n_24));
   AOI21_X1 i_41 (.A(n_116), .B1(n_121), .B2(n_114), .ZN(n_25));
   OAI21_X1 i_42 (.A(n_114), .B1(M[12]), .B2(A[12]), .ZN(n_26));
   NOR2_X1 i_43 (.A1(n_120), .A2(n_111), .ZN(n_27));
   XOR2_X1 i_44 (.A(n_107), .B(n_34), .Z(p_0[16]));
   XOR2_X1 i_45 (.A(n_33), .B(n_30), .Z(p_0[17]));
   XOR2_X1 i_46 (.A(n_31), .B(n_28), .Z(p_0[18]));
   NOR2_X1 i_47 (.A1(n_104), .A2(n_95), .ZN(n_28));
   XNOR2_X1 i_48 (.A(n_35), .B(n_29), .ZN(p_0[19]));
   OAI22_X1 i_49 (.A1(M[18]), .A2(A[18]), .B1(n_95), .B2(n_31), .ZN(n_29));
   AOI21_X1 i_50 (.A(n_105), .B1(M[17]), .B2(A[17]), .ZN(n_30));
   AOI21_X1 i_51 (.A(n_105), .B1(n_99), .B2(n_32), .ZN(n_31));
   INV_X1 i_52 (.A(n_33), .ZN(n_32));
   AOI21_X1 i_53 (.A(n_102), .B1(n_107), .B2(n_100), .ZN(n_33));
   OAI21_X1 i_54 (.A(n_100), .B1(M[16]), .B2(A[16]), .ZN(n_34));
   NOR2_X1 i_55 (.A1(n_106), .A2(n_97), .ZN(n_35));
   XOR2_X1 i_56 (.A(n_93), .B(n_42), .Z(p_0[20]));
   XOR2_X1 i_57 (.A(n_41), .B(n_38), .Z(p_0[21]));
   XOR2_X1 i_58 (.A(n_39), .B(n_36), .Z(p_0[22]));
   NOR2_X1 i_59 (.A1(n_82), .A2(n_72), .ZN(n_36));
   XNOR2_X1 i_60 (.A(n_43), .B(n_37), .ZN(p_0[23]));
   OAI21_X1 i_61 (.A(n_81), .B1(n_72), .B2(n_39), .ZN(n_37));
   NOR2_X1 i_62 (.A1(n_84), .A2(n_74), .ZN(n_38));
   INV_X1 i_63 (.A(n_40), .ZN(n_39));
   OAI21_X1 i_64 (.A(n_83), .B1(n_74), .B2(n_41), .ZN(n_40));
   AOI21_X1 i_65 (.A(n_79), .B1(n_93), .B2(n_76), .ZN(n_41));
   OAI21_X1 i_66 (.A(n_76), .B1(M[20]), .B2(A[20]), .ZN(n_42));
   AOI21_X1 i_67 (.A(n_86), .B1(M[23]), .B2(A[23]), .ZN(n_43));
   XOR2_X1 i_68 (.A(n_51), .B(n_50), .Z(p_0[24]));
   XOR2_X1 i_69 (.A(n_49), .B(n_47), .Z(p_0[25]));
   XNOR2_X1 i_70 (.A(n_45), .B(n_44), .ZN(p_0[26]));
   NOR2_X1 i_71 (.A1(n_91), .A2(n_48), .ZN(n_44));
   OAI21_X1 i_72 (.A(n_66), .B1(M[26]), .B2(A[26]), .ZN(n_45));
   XNOR2_X1 i_73 (.A(n_53), .B(n_46), .ZN(p_0[27]));
   OAI21_X1 i_74 (.A(n_66), .B1(n_90), .B2(n_48), .ZN(n_46));
   AOI21_X1 i_75 (.A(n_91), .B1(M[25]), .B2(A[25]), .ZN(n_47));
   AOI21_X1 i_76 (.A(n_49), .B1(M[25]), .B2(A[25]), .ZN(n_48));
   AOI21_X1 i_77 (.A(n_88), .B1(n_69), .B2(n_51), .ZN(n_49));
   OAI21_X1 i_78 (.A(n_69), .B1(M[24]), .B2(A[24]), .ZN(n_50));
   INV_X1 i_79 (.A(n_52), .ZN(n_51));
   OAI21_X1 i_80 (.A(n_71), .B1(n_93), .B2(n_78), .ZN(n_52));
   OAI22_X1 i_81 (.A1(M[27]), .A2(A[27]), .B1(n_165), .B2(n_162), .ZN(n_53));
   XNOR2_X1 i_82 (.A(n_64), .B(n_63), .ZN(p_0[28]));
   XOR2_X1 i_83 (.A(n_62), .B(n_58), .Z(p_0[29]));
   XNOR2_X1 i_84 (.A(n_55), .B(n_54), .ZN(p_0[30]));
   OAI21_X1 i_85 (.A(n_160), .B1(n_166), .B2(n_163), .ZN(n_54));
   NOR2_X1 i_86 (.A1(n_61), .A2(n_60), .ZN(n_55));
   XOR2_X1 i_87 (.A(n_57), .B(n_56), .Z(p_0[31]));
   XNOR2_X1 i_88 (.A(M[31]), .B(M[30]), .ZN(n_56));
   OAI21_X1 i_89 (.A(n_160), .B1(n_61), .B2(n_59), .ZN(n_57));
   AOI21_X1 i_90 (.A(n_60), .B1(M[29]), .B2(A[29]), .ZN(n_58));
   OAI22_X1 i_91 (.A1(n_166), .A2(n_163), .B1(M[29]), .B2(A[29]), .ZN(n_59));
   NOR2_X1 i_92 (.A1(M[29]), .A2(A[29]), .ZN(n_60));
   AOI21_X1 i_93 (.A(n_62), .B1(M[29]), .B2(A[29]), .ZN(n_61));
   AOI21_X1 i_94 (.A(n_159), .B1(n_64), .B2(n_63), .ZN(n_62));
   AOI21_X1 i_95 (.A(n_159), .B1(M[28]), .B2(A[28]), .ZN(n_63));
   NOR4_X1 i_96 (.A1(n_67), .A2(n_65), .A3(n_70), .A4(n_77), .ZN(n_64));
   OAI22_X1 i_97 (.A1(n_165), .A2(n_162), .B1(n_92), .B2(n_66), .ZN(n_65));
   NAND2_X1 i_98 (.A1(M[26]), .A2(A[26]), .ZN(n_66));
   AOI21_X1 i_99 (.A(n_89), .B1(n_69), .B2(n_68), .ZN(n_67));
   NAND2_X1 i_100 (.A1(M[25]), .A2(A[25]), .ZN(n_68));
   NAND2_X1 i_101 (.A1(M[24]), .A2(A[24]), .ZN(n_69));
   NOR2_X1 i_102 (.A1(n_87), .A2(n_71), .ZN(n_70));
   AOI221_X1 i_103 (.A(n_73), .B1(M[23]), .B2(A[23]), .C1(n_85), .C2(n_72), 
      .ZN(n_71));
   AND2_X1 i_104 (.A1(M[22]), .A2(A[22]), .ZN(n_72));
   AOI21_X1 i_105 (.A(n_80), .B1(n_76), .B2(n_75), .ZN(n_73));
   INV_X1 i_106 (.A(n_75), .ZN(n_74));
   NAND2_X1 i_107 (.A1(M[21]), .A2(A[21]), .ZN(n_75));
   NAND2_X1 i_108 (.A1(M[20]), .A2(A[20]), .ZN(n_76));
   NOR3_X1 i_109 (.A1(n_87), .A2(n_78), .A3(n_93), .ZN(n_77));
   OR2_X1 i_110 (.A1(n_80), .A2(n_79), .ZN(n_78));
   NOR2_X1 i_111 (.A1(M[20]), .A2(A[20]), .ZN(n_79));
   NAND3_X1 i_112 (.A1(n_85), .A2(n_81), .A3(n_83), .ZN(n_80));
   INV_X1 i_113 (.A(n_82), .ZN(n_81));
   NOR2_X1 i_114 (.A1(M[22]), .A2(A[22]), .ZN(n_82));
   INV_X1 i_115 (.A(n_84), .ZN(n_83));
   NOR2_X1 i_116 (.A1(M[21]), .A2(A[21]), .ZN(n_84));
   INV_X1 i_117 (.A(n_86), .ZN(n_85));
   NOR2_X1 i_118 (.A1(M[23]), .A2(A[23]), .ZN(n_86));
   OR2_X1 i_119 (.A1(n_89), .A2(n_88), .ZN(n_87));
   NOR2_X1 i_120 (.A1(M[24]), .A2(A[24]), .ZN(n_88));
   OR2_X1 i_121 (.A1(n_92), .A2(n_90), .ZN(n_89));
   OAI22_X1 i_122 (.A1(M[25]), .A2(A[25]), .B1(M[26]), .B2(A[26]), .ZN(n_90));
   NOR2_X1 i_123 (.A1(M[25]), .A2(A[25]), .ZN(n_91));
   NOR2_X1 i_124 (.A1(M[27]), .A2(A[27]), .ZN(n_92));
   NOR4_X1 i_125 (.A1(n_97), .A2(n_94), .A3(n_98), .A4(n_101), .ZN(n_93));
   NOR2_X1 i_126 (.A1(n_106), .A2(n_96), .ZN(n_94));
   INV_X1 i_127 (.A(n_96), .ZN(n_95));
   NAND2_X1 i_128 (.A1(M[18]), .A2(A[18]), .ZN(n_96));
   AND2_X1 i_129 (.A1(M[19]), .A2(A[19]), .ZN(n_97));
   AOI21_X1 i_130 (.A(n_103), .B1(n_100), .B2(n_99), .ZN(n_98));
   NAND2_X1 i_131 (.A1(M[17]), .A2(A[17]), .ZN(n_99));
   NAND2_X1 i_132 (.A1(M[16]), .A2(A[16]), .ZN(n_100));
   NOR3_X1 i_133 (.A1(n_103), .A2(n_102), .A3(n_107), .ZN(n_101));
   NOR2_X1 i_134 (.A1(M[16]), .A2(A[16]), .ZN(n_102));
   OR3_X1 i_135 (.A1(n_106), .A2(n_104), .A3(n_105), .ZN(n_103));
   NOR2_X1 i_136 (.A1(M[18]), .A2(A[18]), .ZN(n_104));
   NOR2_X1 i_137 (.A1(M[17]), .A2(A[17]), .ZN(n_105));
   NOR2_X1 i_138 (.A1(M[19]), .A2(A[19]), .ZN(n_106));
   NOR4_X1 i_139 (.A1(n_111), .A2(n_108), .A3(n_112), .A4(n_115), .ZN(n_107));
   NOR2_X1 i_140 (.A1(n_120), .A2(n_110), .ZN(n_108));
   INV_X1 i_141 (.A(n_110), .ZN(n_109));
   NAND2_X1 i_142 (.A1(M[14]), .A2(A[14]), .ZN(n_110));
   AND2_X1 i_143 (.A1(M[15]), .A2(A[15]), .ZN(n_111));
   AOI21_X1 i_144 (.A(n_117), .B1(n_114), .B2(n_113), .ZN(n_112));
   NAND2_X1 i_145 (.A1(M[13]), .A2(A[13]), .ZN(n_113));
   NAND2_X1 i_146 (.A1(M[12]), .A2(A[12]), .ZN(n_114));
   NOR3_X1 i_147 (.A1(n_117), .A2(n_116), .A3(n_121), .ZN(n_115));
   NOR2_X1 i_148 (.A1(M[12]), .A2(A[12]), .ZN(n_116));
   OR3_X1 i_149 (.A1(n_120), .A2(n_118), .A3(n_119), .ZN(n_117));
   NOR2_X1 i_150 (.A1(M[14]), .A2(A[14]), .ZN(n_118));
   NOR2_X1 i_151 (.A1(M[13]), .A2(A[13]), .ZN(n_119));
   NOR2_X1 i_152 (.A1(M[15]), .A2(A[15]), .ZN(n_120));
   NOR4_X1 i_153 (.A1(n_125), .A2(n_122), .A3(n_126), .A4(n_129), .ZN(n_121));
   NOR2_X1 i_154 (.A1(n_134), .A2(n_124), .ZN(n_122));
   INV_X1 i_155 (.A(n_124), .ZN(n_123));
   NAND2_X1 i_156 (.A1(M[10]), .A2(A[10]), .ZN(n_124));
   AND2_X1 i_157 (.A1(M[11]), .A2(A[11]), .ZN(n_125));
   AOI21_X1 i_158 (.A(n_131), .B1(n_128), .B2(n_127), .ZN(n_126));
   NAND2_X1 i_159 (.A1(M[9]), .A2(A[9]), .ZN(n_127));
   NAND2_X1 i_160 (.A1(M[8]), .A2(A[8]), .ZN(n_128));
   NOR3_X1 i_161 (.A1(n_131), .A2(n_130), .A3(n_135), .ZN(n_129));
   NOR2_X1 i_162 (.A1(M[8]), .A2(A[8]), .ZN(n_130));
   OR3_X1 i_163 (.A1(n_134), .A2(n_132), .A3(n_133), .ZN(n_131));
   NOR2_X1 i_164 (.A1(M[10]), .A2(A[10]), .ZN(n_132));
   NOR2_X1 i_165 (.A1(M[9]), .A2(A[9]), .ZN(n_133));
   NOR2_X1 i_166 (.A1(M[11]), .A2(A[11]), .ZN(n_134));
   NOR4_X1 i_167 (.A1(n_139), .A2(n_136), .A3(n_140), .A4(n_143), .ZN(n_135));
   NOR2_X1 i_168 (.A1(n_148), .A2(n_138), .ZN(n_136));
   INV_X1 i_169 (.A(n_138), .ZN(n_137));
   NAND2_X1 i_170 (.A1(M[6]), .A2(A[6]), .ZN(n_138));
   AND2_X1 i_171 (.A1(M[7]), .A2(A[7]), .ZN(n_139));
   AOI21_X1 i_172 (.A(n_145), .B1(n_142), .B2(n_141), .ZN(n_140));
   NAND2_X1 i_173 (.A1(M[5]), .A2(A[5]), .ZN(n_141));
   NAND2_X1 i_174 (.A1(M[4]), .A2(A[4]), .ZN(n_142));
   NOR3_X1 i_175 (.A1(n_145), .A2(n_144), .A3(n_149), .ZN(n_143));
   NOR2_X1 i_176 (.A1(M[4]), .A2(A[4]), .ZN(n_144));
   OR3_X1 i_177 (.A1(n_148), .A2(n_146), .A3(n_147), .ZN(n_145));
   NOR2_X1 i_178 (.A1(M[6]), .A2(A[6]), .ZN(n_146));
   NOR2_X1 i_179 (.A1(M[5]), .A2(A[5]), .ZN(n_147));
   NOR2_X1 i_180 (.A1(M[7]), .A2(A[7]), .ZN(n_148));
   NAND2_X1 i_181 (.A1(n_158), .A2(n_150), .ZN(n_149));
   OAI21_X1 i_182 (.A(n_151), .B1(n_164), .B2(n_161), .ZN(n_150));
   OAI22_X1 i_183 (.A1(M[2]), .A2(A[2]), .B1(n_156), .B2(n_152), .ZN(n_151));
   AOI21_X1 i_184 (.A(n_155), .B1(n_154), .B2(n_153), .ZN(n_152));
   NAND2_X1 i_185 (.A1(M[1]), .A2(A[1]), .ZN(n_153));
   NAND2_X1 i_186 (.A1(M[0]), .A2(A[0]), .ZN(n_154));
   NOR2_X1 i_187 (.A1(M[1]), .A2(A[1]), .ZN(n_155));
   INV_X1 i_188 (.A(n_157), .ZN(n_156));
   NAND2_X1 i_189 (.A1(M[2]), .A2(A[2]), .ZN(n_157));
   NAND2_X1 i_190 (.A1(n_164), .A2(n_161), .ZN(n_158));
   NOR2_X1 i_191 (.A1(M[28]), .A2(A[28]), .ZN(n_159));
   NAND2_X1 i_192 (.A1(n_166), .A2(n_163), .ZN(n_160));
   INV_X1 i_193 (.A(A[3]), .ZN(n_161));
   INV_X1 i_194 (.A(A[27]), .ZN(n_162));
   INV_X1 i_195 (.A(A[31]), .ZN(n_163));
   INV_X1 i_196 (.A(M[3]), .ZN(n_164));
   INV_X1 i_197 (.A(M[27]), .ZN(n_165));
   INV_X1 i_198 (.A(M[30]), .ZN(n_166));
endmodule

module Booth(clk, rst, m, q, P);
   input clk;
   input rst;
   input [31:0]m;
   input [31:0]q;
   output [63:0]P;

   wire n_0_0;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_1;
   wire n_0_0_0;
   wire n_0_2;
   wire n_0_0_1;
   wire n_0_3;
   wire n_0_0_2;
   wire n_0_68;
   wire n_0_0_3;
   wire n_0_69;
   wire n_0_0_4;
   wire n_0_70;
   wire n_0_0_5;
   wire n_0_71;
   wire n_0_0_6;
   wire n_0_72;
   wire n_0_0_7;
   wire n_0_73;
   wire n_0_0_8;
   wire n_0_74;
   wire n_0_0_9;
   wire n_0_75;
   wire n_0_0_10;
   wire n_0_76;
   wire n_0_0_11;
   wire n_0_77;
   wire n_0_0_12;
   wire n_0_78;
   wire n_0_0_13;
   wire n_0_79;
   wire n_0_0_14;
   wire n_0_80;
   wire n_0_0_15;
   wire n_0_81;
   wire n_0_0_16;
   wire n_0_82;
   wire n_0_0_17;
   wire n_0_83;
   wire n_0_0_18;
   wire n_0_84;
   wire n_0_0_19;
   wire n_0_85;
   wire n_0_0_20;
   wire n_0_86;
   wire n_0_0_21;
   wire n_0_87;
   wire n_0_0_22;
   wire n_0_88;
   wire n_0_0_23;
   wire n_0_89;
   wire n_0_0_24;
   wire n_0_90;
   wire n_0_0_25;
   wire n_0_91;
   wire n_0_0_26;
   wire n_0_92;
   wire n_0_0_27;
   wire n_0_93;
   wire n_0_0_28;
   wire n_0_94;
   wire n_0_0_29;
   wire n_0_95;
   wire n_0_0_30;
   wire n_0_0_31;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire n_0_130;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire n_0_134;
   wire n_0_135;
   wire n_0_136;
   wire n_0_137;
   wire n_0_138;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_0_32;
   wire n_0_0_33;
   wire n_0_0_34;
   wire n_0_0_35;
   wire n_0_0_36;
   wire n_0_0_37;
   wire n_0_107;
   wire n_0_108;
   wire n_0_0_38;
   wire n_0_109;
   wire n_0_0_39;
   wire n_0_110;
   wire n_0_0_40;
   wire n_0_111;
   wire n_0_0_41;
   wire n_0_112;
   wire n_0_0_42;
   wire n_0_103;
   wire n_0_104;
   wire n_0_0_43;
   wire n_0_0_44;
   wire n_0_0_45;
   wire n_0_0_46;
   wire [31:0]Q;
   wire [31:0]A;
   wire n_0_105;
   wire [31:0]M;
   wire q1;
   wire [5:0]n;
   wire n_0_106;
   wire n_0_113;

   assign P[63] = P[62];

   CLKGATETST_X1 clk_gate_P_reg (.CK(clk), .E(n_0_104), .SE(1'b0), .GCK(n_0_0));
   DFF_X1 \P_reg[63]  (.D(A[31]), .CK(n_0_0), .Q(P[62]), .QN());
   DFF_X1 \P_reg[61]  (.D(A[29]), .CK(n_0_0), .Q(P[61]), .QN());
   DFF_X1 \P_reg[60]  (.D(A[28]), .CK(n_0_0), .Q(P[60]), .QN());
   DFF_X1 \P_reg[59]  (.D(A[27]), .CK(n_0_0), .Q(P[59]), .QN());
   DFF_X1 \P_reg[58]  (.D(A[26]), .CK(n_0_0), .Q(P[58]), .QN());
   DFF_X1 \P_reg[57]  (.D(A[25]), .CK(n_0_0), .Q(P[57]), .QN());
   DFF_X1 \P_reg[56]  (.D(A[24]), .CK(n_0_0), .Q(P[56]), .QN());
   DFF_X1 \P_reg[55]  (.D(A[23]), .CK(n_0_0), .Q(P[55]), .QN());
   DFF_X1 \P_reg[54]  (.D(A[22]), .CK(n_0_0), .Q(P[54]), .QN());
   DFF_X1 \P_reg[53]  (.D(A[21]), .CK(n_0_0), .Q(P[53]), .QN());
   DFF_X1 \P_reg[52]  (.D(A[20]), .CK(n_0_0), .Q(P[52]), .QN());
   DFF_X1 \P_reg[51]  (.D(A[19]), .CK(n_0_0), .Q(P[51]), .QN());
   DFF_X1 \P_reg[50]  (.D(A[18]), .CK(n_0_0), .Q(P[50]), .QN());
   DFF_X1 \P_reg[49]  (.D(A[17]), .CK(n_0_0), .Q(P[49]), .QN());
   DFF_X1 \P_reg[48]  (.D(A[16]), .CK(n_0_0), .Q(P[48]), .QN());
   DFF_X1 \P_reg[47]  (.D(A[15]), .CK(n_0_0), .Q(P[47]), .QN());
   DFF_X1 \P_reg[46]  (.D(A[14]), .CK(n_0_0), .Q(P[46]), .QN());
   DFF_X1 \P_reg[45]  (.D(A[13]), .CK(n_0_0), .Q(P[45]), .QN());
   DFF_X1 \P_reg[44]  (.D(A[12]), .CK(n_0_0), .Q(P[44]), .QN());
   DFF_X1 \P_reg[43]  (.D(A[11]), .CK(n_0_0), .Q(P[43]), .QN());
   DFF_X1 \P_reg[42]  (.D(A[10]), .CK(n_0_0), .Q(P[42]), .QN());
   DFF_X1 \P_reg[41]  (.D(A[9]), .CK(n_0_0), .Q(P[41]), .QN());
   DFF_X1 \P_reg[40]  (.D(A[8]), .CK(n_0_0), .Q(P[40]), .QN());
   DFF_X1 \P_reg[39]  (.D(A[7]), .CK(n_0_0), .Q(P[39]), .QN());
   DFF_X1 \P_reg[38]  (.D(A[6]), .CK(n_0_0), .Q(P[38]), .QN());
   DFF_X1 \P_reg[37]  (.D(A[5]), .CK(n_0_0), .Q(P[37]), .QN());
   DFF_X1 \P_reg[36]  (.D(A[4]), .CK(n_0_0), .Q(P[36]), .QN());
   DFF_X1 \P_reg[35]  (.D(A[3]), .CK(n_0_0), .Q(P[35]), .QN());
   DFF_X1 \P_reg[34]  (.D(A[2]), .CK(n_0_0), .Q(P[34]), .QN());
   DFF_X1 \P_reg[33]  (.D(A[1]), .CK(n_0_0), .Q(P[33]), .QN());
   DFF_X1 \P_reg[32]  (.D(A[0]), .CK(n_0_0), .Q(P[32]), .QN());
   DFF_X1 \P_reg[31]  (.D(Q[31]), .CK(n_0_0), .Q(P[31]), .QN());
   DFF_X1 \P_reg[30]  (.D(Q[30]), .CK(n_0_0), .Q(P[30]), .QN());
   DFF_X1 \P_reg[29]  (.D(Q[29]), .CK(n_0_0), .Q(P[29]), .QN());
   DFF_X1 \P_reg[28]  (.D(Q[28]), .CK(n_0_0), .Q(P[28]), .QN());
   DFF_X1 \P_reg[27]  (.D(Q[27]), .CK(n_0_0), .Q(P[27]), .QN());
   DFF_X1 \P_reg[26]  (.D(Q[26]), .CK(n_0_0), .Q(P[26]), .QN());
   DFF_X1 \P_reg[25]  (.D(Q[25]), .CK(n_0_0), .Q(P[25]), .QN());
   DFF_X1 \P_reg[24]  (.D(Q[24]), .CK(n_0_0), .Q(P[24]), .QN());
   DFF_X1 \P_reg[23]  (.D(Q[23]), .CK(n_0_0), .Q(P[23]), .QN());
   DFF_X1 \P_reg[22]  (.D(Q[22]), .CK(n_0_0), .Q(P[22]), .QN());
   DFF_X1 \P_reg[21]  (.D(Q[21]), .CK(n_0_0), .Q(P[21]), .QN());
   DFF_X1 \P_reg[20]  (.D(Q[20]), .CK(n_0_0), .Q(P[20]), .QN());
   DFF_X1 \P_reg[19]  (.D(Q[19]), .CK(n_0_0), .Q(P[19]), .QN());
   DFF_X1 \P_reg[18]  (.D(Q[18]), .CK(n_0_0), .Q(P[18]), .QN());
   DFF_X1 \P_reg[17]  (.D(Q[17]), .CK(n_0_0), .Q(P[17]), .QN());
   DFF_X1 \P_reg[16]  (.D(Q[16]), .CK(n_0_0), .Q(P[16]), .QN());
   DFF_X1 \P_reg[15]  (.D(Q[15]), .CK(n_0_0), .Q(P[15]), .QN());
   DFF_X1 \P_reg[14]  (.D(Q[14]), .CK(n_0_0), .Q(P[14]), .QN());
   DFF_X1 \P_reg[13]  (.D(Q[13]), .CK(n_0_0), .Q(P[13]), .QN());
   DFF_X1 \P_reg[12]  (.D(Q[12]), .CK(n_0_0), .Q(P[12]), .QN());
   DFF_X1 \P_reg[11]  (.D(Q[11]), .CK(n_0_0), .Q(P[11]), .QN());
   DFF_X1 \P_reg[10]  (.D(Q[10]), .CK(n_0_0), .Q(P[10]), .QN());
   DFF_X1 \P_reg[9]  (.D(Q[9]), .CK(n_0_0), .Q(P[9]), .QN());
   DFF_X1 \P_reg[8]  (.D(Q[8]), .CK(n_0_0), .Q(P[8]), .QN());
   DFF_X1 \P_reg[7]  (.D(Q[7]), .CK(n_0_0), .Q(P[7]), .QN());
   DFF_X1 \P_reg[6]  (.D(Q[6]), .CK(n_0_0), .Q(P[6]), .QN());
   DFF_X1 \P_reg[5]  (.D(Q[5]), .CK(n_0_0), .Q(P[5]), .QN());
   DFF_X1 \P_reg[4]  (.D(Q[4]), .CK(n_0_0), .Q(P[4]), .QN());
   DFF_X1 \P_reg[3]  (.D(Q[3]), .CK(n_0_0), .Q(P[3]), .QN());
   DFF_X1 \P_reg[2]  (.D(Q[2]), .CK(n_0_0), .Q(P[2]), .QN());
   DFF_X1 \P_reg[1]  (.D(Q[1]), .CK(n_0_0), .Q(P[1]), .QN());
   DFF_X1 \P_reg[0]  (.D(Q[0]), .CK(n_0_0), .Q(P[0]), .QN());
   datapath i_0_3 (.A({A[31], uc_0, A[29], A[28], A[27], A[26], A[25], A[24], 
      A[23], A[22], A[21], A[20], A[19], A[18], A[17], A[16], A[15], A[14], 
      A[13], A[12], A[11], A[10], A[9], A[8], A[7], A[6], A[5], A[4], A[3], A[2], 
      A[1], A[0]}), .p_0({n_0_35, n_0_34, n_0_33, n_0_32, n_0_31, n_0_30, n_0_29, 
      n_0_28, n_0_27, n_0_26, n_0_25, n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, 
      n_0_19, n_0_18, n_0_17, n_0_16, n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, 
      n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, n_0_5, n_0_4}), .M(M));
   datapath__0_1 i_0_4 (.M(M), .A({A[31], uc_1, A[29], A[28], A[27], A[26], 
      A[25], A[24], A[23], A[22], A[21], A[20], A[19], A[18], A[17], A[16], 
      A[15], A[14], A[13], A[12], A[11], A[10], A[9], A[8], A[7], A[6], A[5], 
      A[4], A[3], A[2], A[1], A[0]}), .p_0({n_0_67, n_0_66, n_0_65, n_0_64, 
      n_0_63, n_0_62, n_0_61, n_0_60, n_0_59, n_0_58, n_0_57, n_0_56, n_0_55, 
      n_0_54, n_0_53, n_0_52, n_0_51, n_0_50, n_0_49, n_0_48, n_0_47, n_0_46, 
      n_0_45, n_0_44, n_0_43, n_0_42, n_0_41, n_0_40, n_0_39, n_0_38, n_0_37, 
      n_0_36}));
   INV_X1 i_0_0_0 (.A(n_0_0_0), .ZN(n_0_1));
   AOI222_X1 i_0_0_1 (.A1(A[1]), .A2(n_0_0_36), .B1(n_0_0_34), .B2(n_0_37), 
      .C1(n_0_0_33), .C2(n_0_5), .ZN(n_0_0_0));
   INV_X1 i_0_0_2 (.A(n_0_0_1), .ZN(n_0_2));
   AOI222_X1 i_0_0_3 (.A1(A[2]), .A2(n_0_0_36), .B1(n_0_0_34), .B2(n_0_38), 
      .C1(n_0_0_33), .C2(n_0_6), .ZN(n_0_0_1));
   INV_X1 i_0_0_4 (.A(n_0_0_2), .ZN(n_0_3));
   AOI222_X1 i_0_0_5 (.A1(A[3]), .A2(n_0_0_36), .B1(n_0_0_34), .B2(n_0_39), 
      .C1(n_0_0_33), .C2(n_0_7), .ZN(n_0_0_2));
   INV_X1 i_0_0_6 (.A(n_0_0_3), .ZN(n_0_68));
   AOI222_X1 i_0_0_7 (.A1(A[4]), .A2(n_0_0_36), .B1(n_0_0_34), .B2(n_0_40), 
      .C1(n_0_0_33), .C2(n_0_8), .ZN(n_0_0_3));
   INV_X1 i_0_0_8 (.A(n_0_0_4), .ZN(n_0_69));
   AOI222_X1 i_0_0_9 (.A1(A[5]), .A2(n_0_0_36), .B1(n_0_0_34), .B2(n_0_41), 
      .C1(n_0_0_33), .C2(n_0_9), .ZN(n_0_0_4));
   INV_X1 i_0_0_10 (.A(n_0_0_5), .ZN(n_0_70));
   AOI222_X1 i_0_0_11 (.A1(A[6]), .A2(n_0_0_36), .B1(n_0_0_34), .B2(n_0_42), 
      .C1(n_0_0_33), .C2(n_0_10), .ZN(n_0_0_5));
   INV_X1 i_0_0_12 (.A(n_0_0_6), .ZN(n_0_71));
   AOI222_X1 i_0_0_13 (.A1(A[7]), .A2(n_0_0_36), .B1(n_0_0_34), .B2(n_0_43), 
      .C1(n_0_0_33), .C2(n_0_11), .ZN(n_0_0_6));
   INV_X1 i_0_0_14 (.A(n_0_0_7), .ZN(n_0_72));
   AOI222_X1 i_0_0_15 (.A1(A[8]), .A2(n_0_0_36), .B1(n_0_0_34), .B2(n_0_44), 
      .C1(n_0_0_33), .C2(n_0_12), .ZN(n_0_0_7));
   INV_X1 i_0_0_16 (.A(n_0_0_8), .ZN(n_0_73));
   AOI222_X1 i_0_0_17 (.A1(A[9]), .A2(n_0_0_36), .B1(n_0_0_34), .B2(n_0_45), 
      .C1(n_0_0_33), .C2(n_0_13), .ZN(n_0_0_8));
   INV_X1 i_0_0_18 (.A(n_0_0_9), .ZN(n_0_74));
   AOI222_X1 i_0_0_19 (.A1(A[10]), .A2(n_0_0_36), .B1(n_0_0_34), .B2(n_0_46), 
      .C1(n_0_0_33), .C2(n_0_14), .ZN(n_0_0_9));
   INV_X1 i_0_0_20 (.A(n_0_0_10), .ZN(n_0_75));
   AOI222_X1 i_0_0_21 (.A1(A[11]), .A2(n_0_0_36), .B1(n_0_0_34), .B2(n_0_47), 
      .C1(n_0_0_33), .C2(n_0_15), .ZN(n_0_0_10));
   INV_X1 i_0_0_22 (.A(n_0_0_11), .ZN(n_0_76));
   AOI222_X1 i_0_0_23 (.A1(A[12]), .A2(n_0_0_36), .B1(n_0_0_34), .B2(n_0_48), 
      .C1(n_0_0_33), .C2(n_0_16), .ZN(n_0_0_11));
   INV_X1 i_0_0_24 (.A(n_0_0_12), .ZN(n_0_77));
   AOI222_X1 i_0_0_25 (.A1(A[13]), .A2(n_0_0_36), .B1(n_0_0_34), .B2(n_0_49), 
      .C1(n_0_0_33), .C2(n_0_17), .ZN(n_0_0_12));
   INV_X1 i_0_0_26 (.A(n_0_0_13), .ZN(n_0_78));
   AOI222_X1 i_0_0_27 (.A1(A[14]), .A2(n_0_0_36), .B1(n_0_0_34), .B2(n_0_50), 
      .C1(n_0_0_33), .C2(n_0_18), .ZN(n_0_0_13));
   INV_X1 i_0_0_28 (.A(n_0_0_14), .ZN(n_0_79));
   AOI222_X1 i_0_0_29 (.A1(A[15]), .A2(n_0_0_36), .B1(n_0_0_34), .B2(n_0_51), 
      .C1(n_0_0_33), .C2(n_0_19), .ZN(n_0_0_14));
   INV_X1 i_0_0_30 (.A(n_0_0_15), .ZN(n_0_80));
   AOI222_X1 i_0_0_31 (.A1(A[16]), .A2(n_0_0_36), .B1(n_0_0_34), .B2(n_0_52), 
      .C1(n_0_0_33), .C2(n_0_20), .ZN(n_0_0_15));
   INV_X1 i_0_0_32 (.A(n_0_0_16), .ZN(n_0_81));
   AOI222_X1 i_0_0_33 (.A1(A[17]), .A2(n_0_0_36), .B1(n_0_0_34), .B2(n_0_53), 
      .C1(n_0_0_33), .C2(n_0_21), .ZN(n_0_0_16));
   INV_X1 i_0_0_34 (.A(n_0_0_17), .ZN(n_0_82));
   AOI222_X1 i_0_0_35 (.A1(A[18]), .A2(n_0_0_36), .B1(n_0_0_34), .B2(n_0_54), 
      .C1(n_0_0_33), .C2(n_0_22), .ZN(n_0_0_17));
   INV_X1 i_0_0_36 (.A(n_0_0_18), .ZN(n_0_83));
   AOI222_X1 i_0_0_37 (.A1(A[19]), .A2(n_0_0_36), .B1(n_0_0_34), .B2(n_0_55), 
      .C1(n_0_0_33), .C2(n_0_23), .ZN(n_0_0_18));
   INV_X1 i_0_0_38 (.A(n_0_0_19), .ZN(n_0_84));
   AOI222_X1 i_0_0_39 (.A1(A[20]), .A2(n_0_0_36), .B1(n_0_0_34), .B2(n_0_56), 
      .C1(n_0_0_33), .C2(n_0_24), .ZN(n_0_0_19));
   INV_X1 i_0_0_40 (.A(n_0_0_20), .ZN(n_0_85));
   AOI222_X1 i_0_0_41 (.A1(A[21]), .A2(n_0_0_36), .B1(n_0_0_34), .B2(n_0_57), 
      .C1(n_0_0_33), .C2(n_0_25), .ZN(n_0_0_20));
   INV_X1 i_0_0_42 (.A(n_0_0_21), .ZN(n_0_86));
   AOI222_X1 i_0_0_43 (.A1(A[22]), .A2(n_0_0_36), .B1(n_0_0_34), .B2(n_0_58), 
      .C1(n_0_0_33), .C2(n_0_26), .ZN(n_0_0_21));
   INV_X1 i_0_0_44 (.A(n_0_0_22), .ZN(n_0_87));
   AOI222_X1 i_0_0_45 (.A1(A[23]), .A2(n_0_0_36), .B1(n_0_0_34), .B2(n_0_59), 
      .C1(n_0_0_33), .C2(n_0_27), .ZN(n_0_0_22));
   INV_X1 i_0_0_46 (.A(n_0_0_23), .ZN(n_0_88));
   AOI222_X1 i_0_0_47 (.A1(A[24]), .A2(n_0_0_36), .B1(n_0_0_34), .B2(n_0_60), 
      .C1(n_0_0_33), .C2(n_0_28), .ZN(n_0_0_23));
   INV_X1 i_0_0_48 (.A(n_0_0_24), .ZN(n_0_89));
   AOI222_X1 i_0_0_49 (.A1(A[25]), .A2(n_0_0_36), .B1(n_0_0_34), .B2(n_0_61), 
      .C1(n_0_0_33), .C2(n_0_29), .ZN(n_0_0_24));
   INV_X1 i_0_0_50 (.A(n_0_0_25), .ZN(n_0_90));
   AOI222_X1 i_0_0_51 (.A1(A[26]), .A2(n_0_0_36), .B1(n_0_0_34), .B2(n_0_62), 
      .C1(n_0_0_33), .C2(n_0_30), .ZN(n_0_0_25));
   INV_X1 i_0_0_52 (.A(n_0_0_26), .ZN(n_0_91));
   AOI222_X1 i_0_0_53 (.A1(A[27]), .A2(n_0_0_36), .B1(n_0_0_34), .B2(n_0_63), 
      .C1(n_0_0_33), .C2(n_0_31), .ZN(n_0_0_26));
   INV_X1 i_0_0_54 (.A(n_0_0_27), .ZN(n_0_92));
   AOI222_X1 i_0_0_55 (.A1(A[28]), .A2(n_0_0_36), .B1(n_0_0_34), .B2(n_0_64), 
      .C1(n_0_0_33), .C2(n_0_32), .ZN(n_0_0_27));
   INV_X1 i_0_0_56 (.A(n_0_0_28), .ZN(n_0_93));
   AOI222_X1 i_0_0_57 (.A1(A[29]), .A2(n_0_0_36), .B1(n_0_0_34), .B2(n_0_65), 
      .C1(n_0_0_33), .C2(n_0_33), .ZN(n_0_0_28));
   NAND2_X1 i_0_0_58 (.A1(n_0_0_31), .A2(n_0_0_29), .ZN(n_0_94));
   AOI22_X1 i_0_0_59 (.A1(n_0_66), .A2(n_0_0_34), .B1(n_0_0_33), .B2(n_0_34), 
      .ZN(n_0_0_29));
   NAND2_X1 i_0_0_60 (.A1(n_0_0_31), .A2(n_0_0_30), .ZN(n_0_95));
   AOI22_X1 i_0_0_61 (.A1(n_0_67), .A2(n_0_0_34), .B1(n_0_0_33), .B2(n_0_35), 
      .ZN(n_0_0_30));
   NAND2_X1 i_0_0_62 (.A1(A[31]), .A2(n_0_0_36), .ZN(n_0_0_31));
   MUX2_X1 i_0_0_63 (.A(Q[1]), .B(q[0]), .S(rst), .Z(n_0_114));
   MUX2_X1 i_0_0_64 (.A(Q[2]), .B(q[1]), .S(rst), .Z(n_0_115));
   MUX2_X1 i_0_0_65 (.A(Q[3]), .B(q[2]), .S(rst), .Z(n_0_116));
   MUX2_X1 i_0_0_66 (.A(Q[4]), .B(q[3]), .S(rst), .Z(n_0_117));
   MUX2_X1 i_0_0_67 (.A(Q[5]), .B(q[4]), .S(rst), .Z(n_0_118));
   MUX2_X1 i_0_0_68 (.A(Q[6]), .B(q[5]), .S(rst), .Z(n_0_119));
   MUX2_X1 i_0_0_69 (.A(Q[7]), .B(q[6]), .S(rst), .Z(n_0_120));
   MUX2_X1 i_0_0_70 (.A(Q[8]), .B(q[7]), .S(rst), .Z(n_0_121));
   MUX2_X1 i_0_0_71 (.A(Q[9]), .B(q[8]), .S(rst), .Z(n_0_122));
   MUX2_X1 i_0_0_72 (.A(Q[10]), .B(q[9]), .S(rst), .Z(n_0_123));
   MUX2_X1 i_0_0_73 (.A(Q[11]), .B(q[10]), .S(rst), .Z(n_0_124));
   MUX2_X1 i_0_0_74 (.A(Q[12]), .B(q[11]), .S(rst), .Z(n_0_125));
   MUX2_X1 i_0_0_75 (.A(Q[13]), .B(q[12]), .S(rst), .Z(n_0_126));
   MUX2_X1 i_0_0_76 (.A(Q[14]), .B(q[13]), .S(rst), .Z(n_0_127));
   MUX2_X1 i_0_0_77 (.A(Q[15]), .B(q[14]), .S(rst), .Z(n_0_128));
   MUX2_X1 i_0_0_78 (.A(Q[16]), .B(q[15]), .S(rst), .Z(n_0_129));
   MUX2_X1 i_0_0_79 (.A(Q[17]), .B(q[16]), .S(rst), .Z(n_0_130));
   MUX2_X1 i_0_0_80 (.A(Q[18]), .B(q[17]), .S(rst), .Z(n_0_131));
   MUX2_X1 i_0_0_81 (.A(Q[19]), .B(q[18]), .S(rst), .Z(n_0_132));
   MUX2_X1 i_0_0_82 (.A(Q[20]), .B(q[19]), .S(rst), .Z(n_0_133));
   MUX2_X1 i_0_0_83 (.A(Q[21]), .B(q[20]), .S(rst), .Z(n_0_134));
   MUX2_X1 i_0_0_84 (.A(Q[22]), .B(q[21]), .S(rst), .Z(n_0_135));
   MUX2_X1 i_0_0_85 (.A(Q[23]), .B(q[22]), .S(rst), .Z(n_0_136));
   MUX2_X1 i_0_0_86 (.A(Q[24]), .B(q[23]), .S(rst), .Z(n_0_137));
   MUX2_X1 i_0_0_87 (.A(Q[25]), .B(q[24]), .S(rst), .Z(n_0_138));
   MUX2_X1 i_0_0_88 (.A(Q[26]), .B(q[25]), .S(rst), .Z(n_0_96));
   MUX2_X1 i_0_0_89 (.A(Q[27]), .B(q[26]), .S(rst), .Z(n_0_97));
   MUX2_X1 i_0_0_90 (.A(Q[28]), .B(q[27]), .S(rst), .Z(n_0_98));
   MUX2_X1 i_0_0_91 (.A(Q[29]), .B(q[28]), .S(rst), .Z(n_0_99));
   MUX2_X1 i_0_0_92 (.A(Q[30]), .B(q[29]), .S(rst), .Z(n_0_100));
   MUX2_X1 i_0_0_93 (.A(Q[31]), .B(q[30]), .S(rst), .Z(n_0_101));
   NAND2_X1 i_0_0_94 (.A1(n_0_0_32), .A2(n_0_0_35), .ZN(n_0_102));
   AOI222_X1 i_0_0_95 (.A1(rst), .A2(q[31]), .B1(n_0_0_34), .B2(n_0_36), 
      .C1(n_0_0_33), .C2(n_0_4), .ZN(n_0_0_32));
   NOR3_X1 i_0_0_96 (.A1(n_0_0_45), .A2(q1), .A3(rst), .ZN(n_0_0_33));
   NOR3_X1 i_0_0_97 (.A1(n_0_0_46), .A2(Q[0]), .A3(rst), .ZN(n_0_0_34));
   NAND2_X1 i_0_0_98 (.A1(A[0]), .A2(n_0_0_36), .ZN(n_0_0_35));
   NOR2_X1 i_0_0_99 (.A1(n_0_0_37), .A2(rst), .ZN(n_0_0_36));
   XNOR2_X1 i_0_0_100 (.A(n_0_0_46), .B(Q[0]), .ZN(n_0_0_37));
   NOR2_X1 i_0_0_101 (.A1(n[0]), .A2(rst), .ZN(n_0_107));
   NOR2_X1 i_0_0_102 (.A1(rst), .A2(n_0_0_38), .ZN(n_0_108));
   XOR2_X1 i_0_0_103 (.A(n[1]), .B(n[0]), .Z(n_0_0_38));
   AOI21_X1 i_0_0_104 (.A(rst), .B1(n_0_0_44), .B2(n_0_0_39), .ZN(n_0_109));
   OAI21_X1 i_0_0_105 (.A(n[2]), .B1(n[1]), .B2(n[0]), .ZN(n_0_0_39));
   NOR2_X1 i_0_0_106 (.A1(rst), .A2(n_0_0_40), .ZN(n_0_110));
   XOR2_X1 i_0_0_107 (.A(n[3]), .B(n_0_0_44), .Z(n_0_0_40));
   AOI21_X1 i_0_0_108 (.A(rst), .B1(n_0_0_43), .B2(n_0_0_41), .ZN(n_0_111));
   OAI21_X1 i_0_0_109 (.A(n[4]), .B1(n_0_0_44), .B2(n[3]), .ZN(n_0_0_41));
   OAI21_X1 i_0_0_110 (.A(n_0_0_42), .B1(n_0_0_43), .B2(n[5]), .ZN(n_0_112));
   AOI21_X1 i_0_0_111 (.A(rst), .B1(n_0_0_43), .B2(n[5]), .ZN(n_0_0_42));
   NOR2_X1 i_0_0_112 (.A1(n_0_0_45), .A2(rst), .ZN(n_0_103));
   NOR3_X1 i_0_0_113 (.A1(n_0_0_43), .A2(rst), .A3(n[5]), .ZN(n_0_104));
   OR3_X1 i_0_0_114 (.A1(n_0_0_44), .A2(n[3]), .A3(n[4]), .ZN(n_0_0_43));
   OR3_X1 i_0_0_115 (.A1(n[2]), .A2(n[1]), .A3(n[0]), .ZN(n_0_0_44));
   INV_X1 i_0_0_116 (.A(Q[0]), .ZN(n_0_0_45));
   INV_X1 i_0_0_117 (.A(q1), .ZN(n_0_0_46));
   DFF_X1 \Q_reg[31]  (.D(n_0_102), .CK(n_0_106), .Q(Q[31]), .QN());
   DFF_X1 \Q_reg[30]  (.D(n_0_101), .CK(n_0_106), .Q(Q[30]), .QN());
   DFF_X1 \Q_reg[29]  (.D(n_0_100), .CK(n_0_106), .Q(Q[29]), .QN());
   DFF_X1 \Q_reg[28]  (.D(n_0_99), .CK(n_0_106), .Q(Q[28]), .QN());
   DFF_X1 \Q_reg[27]  (.D(n_0_98), .CK(n_0_106), .Q(Q[27]), .QN());
   DFF_X1 \Q_reg[26]  (.D(n_0_97), .CK(n_0_106), .Q(Q[26]), .QN());
   DFF_X1 \Q_reg[25]  (.D(n_0_96), .CK(n_0_106), .Q(Q[25]), .QN());
   DFF_X1 \Q_reg[24]  (.D(n_0_138), .CK(n_0_106), .Q(Q[24]), .QN());
   DFF_X1 \Q_reg[23]  (.D(n_0_137), .CK(n_0_106), .Q(Q[23]), .QN());
   DFF_X1 \Q_reg[22]  (.D(n_0_136), .CK(n_0_106), .Q(Q[22]), .QN());
   DFF_X1 \Q_reg[21]  (.D(n_0_135), .CK(n_0_106), .Q(Q[21]), .QN());
   DFF_X1 \Q_reg[20]  (.D(n_0_134), .CK(n_0_106), .Q(Q[20]), .QN());
   DFF_X1 \Q_reg[19]  (.D(n_0_133), .CK(n_0_106), .Q(Q[19]), .QN());
   DFF_X1 \Q_reg[18]  (.D(n_0_132), .CK(n_0_106), .Q(Q[18]), .QN());
   DFF_X1 \Q_reg[17]  (.D(n_0_131), .CK(n_0_106), .Q(Q[17]), .QN());
   DFF_X1 \Q_reg[16]  (.D(n_0_130), .CK(n_0_106), .Q(Q[16]), .QN());
   DFF_X1 \Q_reg[15]  (.D(n_0_129), .CK(n_0_106), .Q(Q[15]), .QN());
   DFF_X1 \Q_reg[14]  (.D(n_0_128), .CK(n_0_106), .Q(Q[14]), .QN());
   DFF_X1 \Q_reg[13]  (.D(n_0_127), .CK(n_0_106), .Q(Q[13]), .QN());
   DFF_X1 \Q_reg[12]  (.D(n_0_126), .CK(n_0_106), .Q(Q[12]), .QN());
   DFF_X1 \Q_reg[11]  (.D(n_0_125), .CK(n_0_106), .Q(Q[11]), .QN());
   DFF_X1 \Q_reg[10]  (.D(n_0_124), .CK(n_0_106), .Q(Q[10]), .QN());
   DFF_X1 \Q_reg[9]  (.D(n_0_123), .CK(n_0_106), .Q(Q[9]), .QN());
   DFF_X1 \Q_reg[8]  (.D(n_0_122), .CK(n_0_106), .Q(Q[8]), .QN());
   DFF_X1 \Q_reg[7]  (.D(n_0_121), .CK(n_0_106), .Q(Q[7]), .QN());
   DFF_X1 \Q_reg[6]  (.D(n_0_120), .CK(n_0_106), .Q(Q[6]), .QN());
   DFF_X1 \Q_reg[5]  (.D(n_0_119), .CK(n_0_106), .Q(Q[5]), .QN());
   DFF_X1 \Q_reg[4]  (.D(n_0_118), .CK(n_0_106), .Q(Q[4]), .QN());
   DFF_X1 \Q_reg[3]  (.D(n_0_117), .CK(n_0_106), .Q(Q[3]), .QN());
   DFF_X1 \Q_reg[2]  (.D(n_0_116), .CK(n_0_106), .Q(Q[2]), .QN());
   DFF_X1 \Q_reg[1]  (.D(n_0_115), .CK(n_0_106), .Q(Q[1]), .QN());
   DFF_X1 \Q_reg[0]  (.D(n_0_114), .CK(n_0_106), .Q(Q[0]), .QN());
   DFF_X1 \A_reg[31]  (.D(n_0_95), .CK(n_0_106), .Q(A[31]), .QN());
   DFF_X1 \A_reg[29]  (.D(n_0_94), .CK(n_0_106), .Q(A[29]), .QN());
   DFF_X1 \A_reg[28]  (.D(n_0_93), .CK(n_0_106), .Q(A[28]), .QN());
   DFF_X1 \A_reg[27]  (.D(n_0_92), .CK(n_0_106), .Q(A[27]), .QN());
   DFF_X1 \A_reg[26]  (.D(n_0_91), .CK(n_0_106), .Q(A[26]), .QN());
   DFF_X1 \A_reg[25]  (.D(n_0_90), .CK(n_0_106), .Q(A[25]), .QN());
   DFF_X1 \A_reg[24]  (.D(n_0_89), .CK(n_0_106), .Q(A[24]), .QN());
   DFF_X1 \A_reg[23]  (.D(n_0_88), .CK(n_0_106), .Q(A[23]), .QN());
   DFF_X1 \A_reg[22]  (.D(n_0_87), .CK(n_0_106), .Q(A[22]), .QN());
   DFF_X1 \A_reg[21]  (.D(n_0_86), .CK(n_0_106), .Q(A[21]), .QN());
   DFF_X1 \A_reg[20]  (.D(n_0_85), .CK(n_0_106), .Q(A[20]), .QN());
   DFF_X1 \A_reg[19]  (.D(n_0_84), .CK(n_0_106), .Q(A[19]), .QN());
   DFF_X1 \A_reg[18]  (.D(n_0_83), .CK(n_0_106), .Q(A[18]), .QN());
   DFF_X1 \A_reg[17]  (.D(n_0_82), .CK(n_0_106), .Q(A[17]), .QN());
   DFF_X1 \A_reg[16]  (.D(n_0_81), .CK(n_0_106), .Q(A[16]), .QN());
   DFF_X1 \A_reg[15]  (.D(n_0_80), .CK(n_0_106), .Q(A[15]), .QN());
   DFF_X1 \A_reg[14]  (.D(n_0_79), .CK(n_0_106), .Q(A[14]), .QN());
   DFF_X1 \A_reg[13]  (.D(n_0_78), .CK(n_0_106), .Q(A[13]), .QN());
   DFF_X1 \A_reg[12]  (.D(n_0_77), .CK(n_0_106), .Q(A[12]), .QN());
   DFF_X1 \A_reg[11]  (.D(n_0_76), .CK(n_0_106), .Q(A[11]), .QN());
   DFF_X1 \A_reg[10]  (.D(n_0_75), .CK(n_0_106), .Q(A[10]), .QN());
   DFF_X1 \A_reg[9]  (.D(n_0_74), .CK(n_0_106), .Q(A[9]), .QN());
   DFF_X1 \A_reg[8]  (.D(n_0_73), .CK(n_0_106), .Q(A[8]), .QN());
   DFF_X1 \A_reg[7]  (.D(n_0_72), .CK(n_0_106), .Q(A[7]), .QN());
   DFF_X1 \A_reg[6]  (.D(n_0_71), .CK(n_0_106), .Q(A[6]), .QN());
   DFF_X1 \A_reg[5]  (.D(n_0_70), .CK(n_0_106), .Q(A[5]), .QN());
   DFF_X1 \A_reg[4]  (.D(n_0_69), .CK(n_0_106), .Q(A[4]), .QN());
   DFF_X1 \A_reg[3]  (.D(n_0_68), .CK(n_0_106), .Q(A[3]), .QN());
   DFF_X1 \A_reg[2]  (.D(n_0_3), .CK(n_0_106), .Q(A[2]), .QN());
   DFF_X1 \A_reg[1]  (.D(n_0_2), .CK(n_0_106), .Q(A[1]), .QN());
   DFF_X1 \A_reg[0]  (.D(n_0_1), .CK(n_0_106), .Q(A[0]), .QN());
   CLKGATETST_X1 clk_gate_M_reg (.CK(clk), .E(rst), .SE(1'b0), .GCK(n_0_105));
   DFF_X1 \M_reg[31]  (.D(m[31]), .CK(n_0_105), .Q(M[31]), .QN());
   DFF_X1 \M_reg[30]  (.D(m[30]), .CK(n_0_105), .Q(M[30]), .QN());
   DFF_X1 \M_reg[29]  (.D(m[29]), .CK(n_0_105), .Q(M[29]), .QN());
   DFF_X1 \M_reg[28]  (.D(m[28]), .CK(n_0_105), .Q(M[28]), .QN());
   DFF_X1 \M_reg[27]  (.D(m[27]), .CK(n_0_105), .Q(M[27]), .QN());
   DFF_X1 \M_reg[26]  (.D(m[26]), .CK(n_0_105), .Q(M[26]), .QN());
   DFF_X1 \M_reg[25]  (.D(m[25]), .CK(n_0_105), .Q(M[25]), .QN());
   DFF_X1 \M_reg[24]  (.D(m[24]), .CK(n_0_105), .Q(M[24]), .QN());
   DFF_X1 \M_reg[23]  (.D(m[23]), .CK(n_0_105), .Q(M[23]), .QN());
   DFF_X1 \M_reg[22]  (.D(m[22]), .CK(n_0_105), .Q(M[22]), .QN());
   DFF_X1 \M_reg[21]  (.D(m[21]), .CK(n_0_105), .Q(M[21]), .QN());
   DFF_X1 \M_reg[20]  (.D(m[20]), .CK(n_0_105), .Q(M[20]), .QN());
   DFF_X1 \M_reg[19]  (.D(m[19]), .CK(n_0_105), .Q(M[19]), .QN());
   DFF_X1 \M_reg[18]  (.D(m[18]), .CK(n_0_105), .Q(M[18]), .QN());
   DFF_X1 \M_reg[17]  (.D(m[17]), .CK(n_0_105), .Q(M[17]), .QN());
   DFF_X1 \M_reg[16]  (.D(m[16]), .CK(n_0_105), .Q(M[16]), .QN());
   DFF_X1 \M_reg[15]  (.D(m[15]), .CK(n_0_105), .Q(M[15]), .QN());
   DFF_X1 \M_reg[14]  (.D(m[14]), .CK(n_0_105), .Q(M[14]), .QN());
   DFF_X1 \M_reg[13]  (.D(m[13]), .CK(n_0_105), .Q(M[13]), .QN());
   DFF_X1 \M_reg[12]  (.D(m[12]), .CK(n_0_105), .Q(M[12]), .QN());
   DFF_X1 \M_reg[11]  (.D(m[11]), .CK(n_0_105), .Q(M[11]), .QN());
   DFF_X1 \M_reg[10]  (.D(m[10]), .CK(n_0_105), .Q(M[10]), .QN());
   DFF_X1 \M_reg[9]  (.D(m[9]), .CK(n_0_105), .Q(M[9]), .QN());
   DFF_X1 \M_reg[8]  (.D(m[8]), .CK(n_0_105), .Q(M[8]), .QN());
   DFF_X1 \M_reg[7]  (.D(m[7]), .CK(n_0_105), .Q(M[7]), .QN());
   DFF_X1 \M_reg[6]  (.D(m[6]), .CK(n_0_105), .Q(M[6]), .QN());
   DFF_X1 \M_reg[5]  (.D(m[5]), .CK(n_0_105), .Q(M[5]), .QN());
   DFF_X1 \M_reg[4]  (.D(m[4]), .CK(n_0_105), .Q(M[4]), .QN());
   DFF_X1 \M_reg[3]  (.D(m[3]), .CK(n_0_105), .Q(M[3]), .QN());
   DFF_X1 \M_reg[2]  (.D(m[2]), .CK(n_0_105), .Q(M[2]), .QN());
   DFF_X1 \M_reg[1]  (.D(m[1]), .CK(n_0_105), .Q(M[1]), .QN());
   DFF_X1 \M_reg[0]  (.D(m[0]), .CK(n_0_105), .Q(M[0]), .QN());
   DFF_X1 q1_reg (.D(n_0_103), .CK(n_0_106), .Q(q1), .QN());
   DFF_X1 \n_reg[5]  (.D(n_0_112), .CK(n_0_106), .Q(n[5]), .QN());
   DFF_X1 \n_reg[4]  (.D(n_0_111), .CK(n_0_106), .Q(n[4]), .QN());
   DFF_X1 \n_reg[3]  (.D(n_0_110), .CK(n_0_106), .Q(n[3]), .QN());
   DFF_X1 \n_reg[2]  (.D(n_0_109), .CK(n_0_106), .Q(n[2]), .QN());
   DFF_X1 \n_reg[1]  (.D(n_0_108), .CK(n_0_106), .Q(n[1]), .QN());
   DFF_X1 \n_reg[0]  (.D(n_0_107), .CK(n_0_106), .Q(n[0]), .QN());
   CLKGATETST_X1 clk_gate_A_reg (.CK(clk), .E(n_0_113), .SE(1'b0), .GCK(n_0_106));
   INV_X1 i_0_12 (.A(n_0_104), .ZN(n_0_113));
endmodule
