/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Fri Dec 23 16:50:06 2022
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 4250487705 */

module datapath(p_0, op1);
   output [31:0]p_0;
   input [31:0]op1;

   XOR2_X1 i_0 (.A(op1[1]), .B(op1[0]), .Z(p_0[1]));
   AND2_X1 i_1 (.A1(n_29), .A2(n_0), .ZN(p_0[2]));
   OAI21_X1 i_2 (.A(op1[2]), .B1(op1[1]), .B2(op1[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(op1[3]), .B(n_29), .Z(p_0[3]));
   XOR2_X1 i_4 (.A(op1[4]), .B(n_28), .Z(p_0[4]));
   XOR2_X1 i_5 (.A(op1[5]), .B(n_27), .Z(p_0[5]));
   AND2_X1 i_6 (.A1(n_26), .A2(n_1), .ZN(p_0[6]));
   OAI21_X1 i_7 (.A(op1[6]), .B1(n_27), .B2(op1[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(op1[7]), .B(n_26), .Z(p_0[7]));
   XOR2_X1 i_9 (.A(op1[8]), .B(n_25), .Z(p_0[8]));
   AND2_X1 i_10 (.A1(n_24), .A2(n_2), .ZN(p_0[9]));
   OAI21_X1 i_11 (.A(op1[9]), .B1(n_25), .B2(op1[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(op1[10]), .B(n_24), .Z(p_0[10]));
   XNOR2_X1 i_13 (.A(op1[11]), .B(n_23), .ZN(p_0[11]));
   XOR2_X1 i_14 (.A(op1[12]), .B(n_22), .Z(p_0[12]));
   XNOR2_X1 i_15 (.A(op1[13]), .B(n_21), .ZN(p_0[13]));
   XNOR2_X1 i_16 (.A(op1[14]), .B(n_20), .ZN(p_0[14]));
   XOR2_X1 i_17 (.A(op1[15]), .B(n_19), .Z(p_0[15]));
   AND2_X1 i_18 (.A1(n_18), .A2(n_3), .ZN(p_0[16]));
   OAI21_X1 i_19 (.A(op1[16]), .B1(n_19), .B2(op1[15]), .ZN(n_3));
   XOR2_X1 i_20 (.A(op1[17]), .B(n_18), .Z(p_0[17]));
   XOR2_X1 i_21 (.A(op1[18]), .B(n_17), .Z(p_0[18]));
   XNOR2_X1 i_22 (.A(op1[19]), .B(n_16), .ZN(p_0[19]));
   XNOR2_X1 i_23 (.A(op1[20]), .B(n_15), .ZN(p_0[20]));
   XNOR2_X1 i_24 (.A(op1[21]), .B(n_14), .ZN(p_0[21]));
   XOR2_X1 i_25 (.A(op1[22]), .B(n_13), .Z(p_0[22]));
   XOR2_X1 i_26 (.A(op1[23]), .B(n_12), .Z(p_0[23]));
   XNOR2_X1 i_27 (.A(op1[24]), .B(n_11), .ZN(p_0[24]));
   XNOR2_X1 i_28 (.A(op1[25]), .B(n_10), .ZN(p_0[25]));
   XOR2_X1 i_29 (.A(op1[26]), .B(n_9), .Z(p_0[26]));
   AND2_X1 i_30 (.A1(n_8), .A2(n_4), .ZN(p_0[27]));
   OAI21_X1 i_31 (.A(op1[27]), .B1(n_9), .B2(op1[26]), .ZN(n_4));
   XOR2_X1 i_32 (.A(op1[28]), .B(n_8), .Z(p_0[28]));
   XNOR2_X1 i_33 (.A(op1[29]), .B(n_7), .ZN(p_0[29]));
   XNOR2_X1 i_34 (.A(op1[30]), .B(n_6), .ZN(p_0[30]));
   XNOR2_X1 i_35 (.A(op1[31]), .B(n_5), .ZN(p_0[31]));
   NOR4_X1 i_36 (.A1(n_8), .A2(op1[28]), .A3(op1[29]), .A4(op1[30]), .ZN(n_5));
   NOR3_X1 i_37 (.A1(n_8), .A2(op1[28]), .A3(op1[29]), .ZN(n_6));
   NOR2_X1 i_38 (.A1(n_8), .A2(op1[28]), .ZN(n_7));
   OR3_X1 i_39 (.A1(n_9), .A2(op1[26]), .A3(op1[27]), .ZN(n_8));
   NAND2_X1 i_40 (.A1(n_10), .A2(n_33), .ZN(n_9));
   NOR3_X1 i_41 (.A1(n_12), .A2(op1[23]), .A3(op1[24]), .ZN(n_10));
   NOR2_X1 i_42 (.A1(n_12), .A2(op1[23]), .ZN(n_11));
   OR2_X1 i_43 (.A1(n_13), .A2(op1[22]), .ZN(n_12));
   NAND2_X1 i_44 (.A1(n_14), .A2(n_32), .ZN(n_13));
   NOR4_X1 i_45 (.A1(n_17), .A2(op1[18]), .A3(op1[19]), .A4(op1[20]), .ZN(n_14));
   NOR3_X1 i_46 (.A1(n_17), .A2(op1[18]), .A3(op1[19]), .ZN(n_15));
   NOR2_X1 i_47 (.A1(n_17), .A2(op1[18]), .ZN(n_16));
   OR2_X1 i_48 (.A1(n_18), .A2(op1[17]), .ZN(n_17));
   OR3_X1 i_49 (.A1(n_19), .A2(op1[15]), .A3(op1[16]), .ZN(n_18));
   NAND2_X1 i_50 (.A1(n_20), .A2(n_31), .ZN(n_19));
   NOR3_X1 i_51 (.A1(n_22), .A2(op1[12]), .A3(op1[13]), .ZN(n_20));
   NOR2_X1 i_52 (.A1(n_22), .A2(op1[12]), .ZN(n_21));
   NAND2_X1 i_53 (.A1(n_23), .A2(n_30), .ZN(n_22));
   NOR2_X1 i_54 (.A1(n_24), .A2(op1[10]), .ZN(n_23));
   OR3_X1 i_55 (.A1(n_25), .A2(op1[8]), .A3(op1[9]), .ZN(n_24));
   OR2_X1 i_56 (.A1(n_26), .A2(op1[7]), .ZN(n_25));
   OR3_X1 i_57 (.A1(n_27), .A2(op1[5]), .A3(op1[6]), .ZN(n_26));
   OR2_X1 i_58 (.A1(n_28), .A2(op1[4]), .ZN(n_27));
   OR2_X1 i_59 (.A1(n_29), .A2(op1[3]), .ZN(n_28));
   OR3_X1 i_60 (.A1(op1[2]), .A2(op1[1]), .A3(op1[0]), .ZN(n_29));
   INV_X1 i_61 (.A(op1[11]), .ZN(n_30));
   INV_X1 i_62 (.A(op1[14]), .ZN(n_31));
   INV_X1 i_63 (.A(op1[21]), .ZN(n_32));
   INV_X1 i_64 (.A(op1[25]), .ZN(n_33));
endmodule

module datapath__0_16(p_0, adder, p_1);
   input [63:0]p_0;
   input [63:0]adder;
   output [63:0]p_1;

   INV_X1 i_0 (.A(n_0), .ZN(p_1[0]));
   OAI21_X1 i_1 (.A(n_367), .B1(p_0[0]), .B2(adder[0]), .ZN(n_0));
   XOR2_X1 i_2 (.A(n_367), .B(n_1), .Z(p_1[1]));
   OAI21_X1 i_3 (.A(n_366), .B1(p_0[1]), .B2(adder[1]), .ZN(n_1));
   XNOR2_X1 i_4 (.A(n_365), .B(n_2), .ZN(p_1[2]));
   OAI21_X1 i_5 (.A(n_370), .B1(p_0[2]), .B2(adder[2]), .ZN(n_2));
   XOR2_X1 i_6 (.A(n_364), .B(n_3), .Z(p_1[3]));
   OAI21_X1 i_7 (.A(n_371), .B1(n_376), .B2(n_373), .ZN(n_3));
   XOR2_X1 i_8 (.A(n_362), .B(n_10), .Z(p_1[4]));
   XOR2_X1 i_9 (.A(n_9), .B(n_6), .Z(p_1[5]));
   XOR2_X1 i_10 (.A(n_7), .B(n_4), .Z(p_1[6]));
   NOR2_X1 i_11 (.A1(n_359), .A2(n_350), .ZN(n_4));
   XNOR2_X1 i_12 (.A(n_11), .B(n_5), .ZN(p_1[7]));
   OAI22_X1 i_13 (.A1(p_0[6]), .A2(adder[6]), .B1(n_350), .B2(n_7), .ZN(n_5));
   AOI21_X1 i_14 (.A(n_360), .B1(p_0[5]), .B2(adder[5]), .ZN(n_6));
   AOI21_X1 i_15 (.A(n_360), .B1(n_354), .B2(n_8), .ZN(n_7));
   INV_X1 i_16 (.A(n_9), .ZN(n_8));
   AOI21_X1 i_17 (.A(n_357), .B1(n_362), .B2(n_355), .ZN(n_9));
   OAI21_X1 i_18 (.A(n_355), .B1(p_0[4]), .B2(adder[4]), .ZN(n_10));
   NOR2_X1 i_19 (.A1(n_361), .A2(n_352), .ZN(n_11));
   XNOR2_X1 i_20 (.A(n_348), .B(n_18), .ZN(p_1[8]));
   XOR2_X1 i_21 (.A(n_17), .B(n_14), .Z(p_1[9]));
   XOR2_X1 i_22 (.A(n_15), .B(n_12), .Z(p_1[10]));
   NOR2_X1 i_23 (.A1(n_345), .A2(n_336), .ZN(n_12));
   XNOR2_X1 i_24 (.A(n_19), .B(n_13), .ZN(p_1[11]));
   OAI22_X1 i_25 (.A1(p_0[10]), .A2(adder[10]), .B1(n_336), .B2(n_15), .ZN(n_13));
   AOI21_X1 i_26 (.A(n_346), .B1(p_0[9]), .B2(adder[9]), .ZN(n_14));
   AOI21_X1 i_27 (.A(n_346), .B1(n_340), .B2(n_16), .ZN(n_15));
   INV_X1 i_28 (.A(n_17), .ZN(n_16));
   AOI21_X1 i_29 (.A(n_343), .B1(n_348), .B2(n_341), .ZN(n_17));
   AOI21_X1 i_30 (.A(n_343), .B1(p_0[8]), .B2(adder[8]), .ZN(n_18));
   NOR2_X1 i_31 (.A1(n_347), .A2(n_338), .ZN(n_19));
   XOR2_X1 i_32 (.A(n_334), .B(n_26), .Z(p_1[12]));
   XOR2_X1 i_33 (.A(n_25), .B(n_22), .Z(p_1[13]));
   XOR2_X1 i_34 (.A(n_23), .B(n_20), .Z(p_1[14]));
   NOR2_X1 i_35 (.A1(n_331), .A2(n_322), .ZN(n_20));
   XNOR2_X1 i_36 (.A(n_27), .B(n_21), .ZN(p_1[15]));
   OAI22_X1 i_37 (.A1(p_0[14]), .A2(adder[14]), .B1(n_322), .B2(n_23), .ZN(n_21));
   AOI21_X1 i_38 (.A(n_332), .B1(p_0[13]), .B2(adder[13]), .ZN(n_22));
   AOI21_X1 i_39 (.A(n_332), .B1(n_326), .B2(n_24), .ZN(n_23));
   INV_X1 i_40 (.A(n_25), .ZN(n_24));
   AOI21_X1 i_41 (.A(n_329), .B1(n_334), .B2(n_327), .ZN(n_25));
   OAI21_X1 i_42 (.A(n_327), .B1(p_0[12]), .B2(adder[12]), .ZN(n_26));
   NOR2_X1 i_43 (.A1(n_333), .A2(n_324), .ZN(n_27));
   XOR2_X1 i_44 (.A(n_320), .B(n_34), .Z(p_1[16]));
   XOR2_X1 i_45 (.A(n_33), .B(n_30), .Z(p_1[17]));
   XOR2_X1 i_46 (.A(n_31), .B(n_28), .Z(p_1[18]));
   NOR2_X1 i_47 (.A1(n_286), .A2(n_276), .ZN(n_28));
   XNOR2_X1 i_48 (.A(n_35), .B(n_29), .ZN(p_1[19]));
   OAI21_X1 i_49 (.A(n_285), .B1(n_276), .B2(n_31), .ZN(n_29));
   NOR2_X1 i_50 (.A1(n_288), .A2(n_278), .ZN(n_30));
   INV_X1 i_51 (.A(n_32), .ZN(n_31));
   OAI21_X1 i_52 (.A(n_287), .B1(n_278), .B2(n_33), .ZN(n_32));
   AOI21_X1 i_53 (.A(n_283), .B1(n_320), .B2(n_280), .ZN(n_33));
   OAI21_X1 i_54 (.A(n_280), .B1(p_0[16]), .B2(adder[16]), .ZN(n_34));
   AOI21_X1 i_55 (.A(n_290), .B1(p_0[19]), .B2(adder[19]), .ZN(n_35));
   XOR2_X1 i_56 (.A(n_63), .B(n_42), .Z(p_1[20]));
   XOR2_X1 i_57 (.A(n_41), .B(n_38), .Z(p_1[21]));
   XOR2_X1 i_58 (.A(n_39), .B(n_36), .Z(p_1[22]));
   NOR2_X1 i_59 (.A1(n_314), .A2(n_258), .ZN(n_36));
   XNOR2_X1 i_60 (.A(n_43), .B(n_37), .ZN(p_1[23]));
   OAI21_X1 i_61 (.A(n_313), .B1(n_258), .B2(n_39), .ZN(n_37));
   NOR2_X1 i_62 (.A1(n_316), .A2(n_260), .ZN(n_38));
   INV_X1 i_63 (.A(n_40), .ZN(n_39));
   OAI21_X1 i_64 (.A(n_315), .B1(n_260), .B2(n_41), .ZN(n_40));
   AOI21_X1 i_65 (.A(n_319), .B1(n_262), .B2(n_63), .ZN(n_41));
   OAI21_X1 i_66 (.A(n_262), .B1(p_0[20]), .B2(adder[20]), .ZN(n_42));
   AOI21_X1 i_67 (.A(n_318), .B1(p_0[23]), .B2(adder[23]), .ZN(n_43));
   XOR2_X1 i_68 (.A(n_61), .B(n_50), .Z(p_1[24]));
   XOR2_X1 i_69 (.A(n_49), .B(n_46), .Z(p_1[25]));
   XOR2_X1 i_70 (.A(n_47), .B(n_44), .Z(p_1[26]));
   NOR2_X1 i_71 (.A1(n_297), .A2(n_270), .ZN(n_44));
   XNOR2_X1 i_72 (.A(n_51), .B(n_45), .ZN(p_1[27]));
   OAI21_X1 i_73 (.A(n_296), .B1(n_270), .B2(n_47), .ZN(n_45));
   NOR2_X1 i_74 (.A1(n_299), .A2(n_272), .ZN(n_46));
   INV_X1 i_75 (.A(n_48), .ZN(n_47));
   OAI21_X1 i_76 (.A(n_298), .B1(n_272), .B2(n_49), .ZN(n_48));
   AOI21_X1 i_77 (.A(n_294), .B1(n_274), .B2(n_61), .ZN(n_49));
   OAI21_X1 i_78 (.A(n_274), .B1(p_0[24]), .B2(adder[24]), .ZN(n_50));
   AOI21_X1 i_79 (.A(n_301), .B1(p_0[27]), .B2(adder[27]), .ZN(n_51));
   XOR2_X1 i_80 (.A(n_59), .B(n_58), .Z(p_1[28]));
   XOR2_X1 i_81 (.A(n_57), .B(n_54), .Z(p_1[29]));
   XOR2_X1 i_82 (.A(n_55), .B(n_52), .Z(p_1[30]));
   NOR2_X1 i_83 (.A1(n_306), .A2(n_264), .ZN(n_52));
   XOR2_X1 i_84 (.A(n_65), .B(n_53), .Z(p_1[31]));
   OAI21_X1 i_85 (.A(n_305), .B1(n_264), .B2(n_55), .ZN(n_53));
   NOR2_X1 i_86 (.A1(n_308), .A2(n_267), .ZN(n_54));
   INV_X1 i_87 (.A(n_56), .ZN(n_55));
   OAI21_X1 i_88 (.A(n_307), .B1(n_267), .B2(n_57), .ZN(n_56));
   AOI21_X1 i_89 (.A(n_303), .B1(n_268), .B2(n_59), .ZN(n_57));
   OAI21_X1 i_90 (.A(n_268), .B1(p_0[28]), .B2(adder[28]), .ZN(n_58));
   INV_X1 i_91 (.A(n_60), .ZN(n_59));
   OAI21_X1 i_92 (.A(n_269), .B1(n_293), .B2(n_61), .ZN(n_60));
   INV_X1 i_93 (.A(n_62), .ZN(n_61));
   OAI21_X1 i_94 (.A(n_257), .B1(n_311), .B2(n_63), .ZN(n_62));
   INV_X1 i_95 (.A(n_64), .ZN(n_63));
   OAI21_X1 i_96 (.A(n_275), .B1(n_320), .B2(n_282), .ZN(n_64));
   OAI21_X1 i_97 (.A(n_309), .B1(n_377), .B2(n_374), .ZN(n_65));
   XOR2_X1 i_98 (.A(n_255), .B(n_72), .Z(p_1[32]));
   XOR2_X1 i_99 (.A(n_71), .B(n_68), .Z(p_1[33]));
   XOR2_X1 i_100 (.A(n_69), .B(n_66), .Z(p_1[34]));
   NOR2_X1 i_101 (.A1(n_224), .A2(n_214), .ZN(n_66));
   XNOR2_X1 i_102 (.A(n_73), .B(n_67), .ZN(p_1[35]));
   OAI21_X1 i_103 (.A(n_223), .B1(n_214), .B2(n_69), .ZN(n_67));
   NOR2_X1 i_104 (.A1(n_226), .A2(n_216), .ZN(n_68));
   INV_X1 i_105 (.A(n_70), .ZN(n_69));
   OAI21_X1 i_106 (.A(n_225), .B1(n_216), .B2(n_71), .ZN(n_70));
   AOI21_X1 i_107 (.A(n_221), .B1(n_255), .B2(n_218), .ZN(n_71));
   OAI21_X1 i_108 (.A(n_218), .B1(p_0[32]), .B2(adder[32]), .ZN(n_72));
   AOI21_X1 i_109 (.A(n_228), .B1(p_0[35]), .B2(adder[35]), .ZN(n_73));
   XOR2_X1 i_110 (.A(n_101), .B(n_80), .Z(p_1[36]));
   XOR2_X1 i_111 (.A(n_79), .B(n_76), .Z(p_1[37]));
   XOR2_X1 i_112 (.A(n_77), .B(n_74), .Z(p_1[38]));
   NOR2_X1 i_113 (.A1(n_249), .A2(n_207), .ZN(n_74));
   XNOR2_X1 i_114 (.A(n_81), .B(n_75), .ZN(p_1[39]));
   OAI21_X1 i_115 (.A(n_248), .B1(n_207), .B2(n_77), .ZN(n_75));
   NOR2_X1 i_116 (.A1(n_251), .A2(n_209), .ZN(n_76));
   INV_X1 i_117 (.A(n_78), .ZN(n_77));
   OAI21_X1 i_118 (.A(n_250), .B1(n_209), .B2(n_79), .ZN(n_78));
   AOI21_X1 i_119 (.A(n_254), .B1(n_211), .B2(n_101), .ZN(n_79));
   OAI21_X1 i_120 (.A(n_211), .B1(p_0[36]), .B2(adder[36]), .ZN(n_80));
   AOI21_X1 i_121 (.A(n_253), .B1(p_0[39]), .B2(adder[39]), .ZN(n_81));
   XOR2_X1 i_122 (.A(n_99), .B(n_88), .Z(p_1[40]));
   XOR2_X1 i_123 (.A(n_87), .B(n_84), .Z(p_1[41]));
   XOR2_X1 i_124 (.A(n_85), .B(n_82), .Z(p_1[42]));
   NOR2_X1 i_125 (.A1(n_235), .A2(n_193), .ZN(n_82));
   XNOR2_X1 i_126 (.A(n_89), .B(n_83), .ZN(p_1[43]));
   OAI21_X1 i_127 (.A(n_234), .B1(n_193), .B2(n_85), .ZN(n_83));
   NOR2_X1 i_128 (.A1(n_237), .A2(n_195), .ZN(n_84));
   INV_X1 i_129 (.A(n_86), .ZN(n_85));
   OAI21_X1 i_130 (.A(n_236), .B1(n_195), .B2(n_87), .ZN(n_86));
   AOI21_X1 i_131 (.A(n_232), .B1(n_197), .B2(n_99), .ZN(n_87));
   OAI21_X1 i_132 (.A(n_197), .B1(p_0[40]), .B2(adder[40]), .ZN(n_88));
   AOI21_X1 i_133 (.A(n_239), .B1(p_0[43]), .B2(adder[43]), .ZN(n_89));
   XNOR2_X1 i_134 (.A(n_98), .B(n_97), .ZN(p_1[44]));
   XOR2_X1 i_135 (.A(n_95), .B(n_94), .Z(p_1[45]));
   XNOR2_X1 i_136 (.A(n_91), .B(n_90), .ZN(p_1[46]));
   OAI22_X1 i_137 (.A1(p_0[45]), .A2(adder[45]), .B1(n_203), .B2(n_95), .ZN(n_90));
   NOR2_X1 i_138 (.A1(n_243), .A2(n_200), .ZN(n_91));
   XNOR2_X1 i_139 (.A(n_103), .B(n_92), .ZN(p_1[47]));
   OAI21_X1 i_140 (.A(n_93), .B1(n_242), .B2(n_200), .ZN(n_92));
   NAND3_X1 i_141 (.A1(n_201), .A2(n_94), .A3(n_96), .ZN(n_93));
   NOR2_X1 i_142 (.A1(n_244), .A2(n_203), .ZN(n_94));
   INV_X1 i_143 (.A(n_96), .ZN(n_95));
   OAI22_X1 i_144 (.A1(p_0[44]), .A2(adder[44]), .B1(n_204), .B2(n_98), .ZN(n_96));
   OAI21_X1 i_145 (.A(n_205), .B1(p_0[44]), .B2(adder[44]), .ZN(n_97));
   OAI21_X1 i_146 (.A(n_192), .B1(n_231), .B2(n_99), .ZN(n_98));
   INV_X1 i_147 (.A(n_100), .ZN(n_99));
   OAI21_X1 i_148 (.A(n_206), .B1(n_246), .B2(n_101), .ZN(n_100));
   INV_X1 i_149 (.A(n_102), .ZN(n_101));
   OAI21_X1 i_150 (.A(n_213), .B1(n_255), .B2(n_220), .ZN(n_102));
   AOI21_X1 i_151 (.A(n_245), .B1(p_0[47]), .B2(adder[47]), .ZN(n_103));
   XOR2_X1 i_152 (.A(n_190), .B(n_110), .Z(p_1[48]));
   XOR2_X1 i_153 (.A(n_109), .B(n_106), .Z(p_1[49]));
   XOR2_X1 i_154 (.A(n_107), .B(n_104), .Z(p_1[50]));
   NOR2_X1 i_155 (.A1(n_187), .A2(n_178), .ZN(n_104));
   XNOR2_X1 i_156 (.A(n_111), .B(n_105), .ZN(p_1[51]));
   OAI22_X1 i_157 (.A1(p_0[50]), .A2(adder[50]), .B1(n_178), .B2(n_107), 
      .ZN(n_105));
   AOI21_X1 i_158 (.A(n_188), .B1(p_0[49]), .B2(adder[49]), .ZN(n_106));
   AOI21_X1 i_159 (.A(n_188), .B1(n_182), .B2(n_108), .ZN(n_107));
   INV_X1 i_160 (.A(n_109), .ZN(n_108));
   AOI21_X1 i_161 (.A(n_185), .B1(n_190), .B2(n_183), .ZN(n_109));
   OAI21_X1 i_162 (.A(n_183), .B1(p_0[48]), .B2(adder[48]), .ZN(n_110));
   NOR2_X1 i_163 (.A1(n_189), .A2(n_180), .ZN(n_111));
   XOR2_X1 i_164 (.A(n_176), .B(n_118), .Z(p_1[52]));
   XOR2_X1 i_165 (.A(n_117), .B(n_114), .Z(p_1[53]));
   XOR2_X1 i_166 (.A(n_115), .B(n_112), .Z(p_1[54]));
   NOR2_X1 i_167 (.A1(n_165), .A2(n_155), .ZN(n_112));
   XNOR2_X1 i_168 (.A(n_119), .B(n_113), .ZN(p_1[55]));
   OAI21_X1 i_169 (.A(n_164), .B1(n_155), .B2(n_115), .ZN(n_113));
   NOR2_X1 i_170 (.A1(n_167), .A2(n_157), .ZN(n_114));
   INV_X1 i_171 (.A(n_116), .ZN(n_115));
   OAI21_X1 i_172 (.A(n_166), .B1(n_157), .B2(n_117), .ZN(n_116));
   AOI21_X1 i_173 (.A(n_162), .B1(n_176), .B2(n_159), .ZN(n_117));
   OAI21_X1 i_174 (.A(n_159), .B1(p_0[52]), .B2(adder[52]), .ZN(n_118));
   AOI21_X1 i_175 (.A(n_169), .B1(p_0[55]), .B2(adder[55]), .ZN(n_119));
   XNOR2_X1 i_176 (.A(n_128), .B(n_127), .ZN(p_1[56]));
   XOR2_X1 i_177 (.A(n_125), .B(n_124), .Z(p_1[57]));
   XNOR2_X1 i_178 (.A(n_121), .B(n_120), .ZN(p_1[58]));
   OAI22_X1 i_179 (.A1(p_0[57]), .A2(adder[57]), .B1(n_150), .B2(n_125), 
      .ZN(n_120));
   NOR2_X1 i_180 (.A1(n_173), .A2(n_146), .ZN(n_121));
   XNOR2_X1 i_181 (.A(n_129), .B(n_122), .ZN(p_1[59]));
   OAI21_X1 i_182 (.A(n_123), .B1(n_172), .B2(n_146), .ZN(n_122));
   NAND3_X1 i_183 (.A1(n_147), .A2(n_124), .A3(n_126), .ZN(n_123));
   NOR2_X1 i_184 (.A1(n_174), .A2(n_150), .ZN(n_124));
   INV_X1 i_185 (.A(n_126), .ZN(n_125));
   OAI22_X1 i_186 (.A1(p_0[56]), .A2(adder[56]), .B1(n_151), .B2(n_128), 
      .ZN(n_126));
   OAI21_X1 i_187 (.A(n_152), .B1(p_0[56]), .B2(adder[56]), .ZN(n_127));
   OAI21_X1 i_188 (.A(n_154), .B1(n_176), .B2(n_161), .ZN(n_128));
   AOI21_X1 i_189 (.A(n_175), .B1(p_0[59]), .B2(adder[59]), .ZN(n_129));
   XNOR2_X1 i_190 (.A(n_144), .B(n_143), .ZN(p_1[60]));
   AOI22_X1 i_191 (.A1(n_141), .A2(n_136), .B1(n_142), .B2(n_137), .ZN(p_1[61]));
   XNOR2_X1 i_192 (.A(n_131), .B(n_130), .ZN(p_1[62]));
   AOI22_X1 i_193 (.A1(p_0[61]), .A2(adder[61]), .B1(n_142), .B2(n_138), 
      .ZN(n_130));
   AOI21_X1 i_194 (.A(n_140), .B1(p_0[61]), .B2(adder[62]), .ZN(n_131));
   XNOR2_X1 i_195 (.A(n_133), .B(n_132), .ZN(p_1[63]));
   XOR2_X1 i_196 (.A(adder[63]), .B(adder[62]), .Z(n_132));
   AOI221_X1 i_197 (.A(n_134), .B1(p_0[61]), .B2(adder[62]), .C1(n_141), 
      .C2(n_135), .ZN(n_133));
   NOR2_X1 i_198 (.A1(n_140), .A2(n_138), .ZN(n_134));
   NOR2_X1 i_199 (.A1(n_140), .A2(n_136), .ZN(n_135));
   INV_X1 i_200 (.A(n_137), .ZN(n_136));
   AOI21_X1 i_201 (.A(n_139), .B1(p_0[61]), .B2(adder[61]), .ZN(n_137));
   INV_X1 i_202 (.A(n_139), .ZN(n_138));
   NOR2_X1 i_203 (.A1(p_0[61]), .A2(adder[61]), .ZN(n_139));
   NOR2_X1 i_204 (.A1(p_0[61]), .A2(adder[62]), .ZN(n_140));
   INV_X1 i_205 (.A(n_142), .ZN(n_141));
   AOI21_X1 i_206 (.A(n_372), .B1(n_144), .B2(n_143), .ZN(n_142));
   AOI21_X1 i_207 (.A(n_372), .B1(p_0[60]), .B2(adder[60]), .ZN(n_143));
   NOR4_X1 i_208 (.A1(n_148), .A2(n_145), .A3(n_153), .A4(n_160), .ZN(n_144));
   OAI22_X1 i_209 (.A1(n_378), .A2(n_375), .B1(n_175), .B2(n_147), .ZN(n_145));
   INV_X1 i_210 (.A(n_147), .ZN(n_146));
   NAND2_X1 i_211 (.A1(p_0[58]), .A2(adder[58]), .ZN(n_147));
   INV_X1 i_212 (.A(n_149), .ZN(n_148));
   OAI21_X1 i_213 (.A(n_171), .B1(n_151), .B2(n_150), .ZN(n_149));
   AND2_X1 i_214 (.A1(p_0[57]), .A2(adder[57]), .ZN(n_150));
   INV_X1 i_215 (.A(n_152), .ZN(n_151));
   NAND2_X1 i_216 (.A1(p_0[56]), .A2(adder[56]), .ZN(n_152));
   NOR2_X1 i_217 (.A1(n_170), .A2(n_154), .ZN(n_153));
   AOI221_X1 i_218 (.A(n_156), .B1(p_0[55]), .B2(adder[55]), .C1(n_168), 
      .C2(n_155), .ZN(n_154));
   AND2_X1 i_219 (.A1(p_0[54]), .A2(adder[54]), .ZN(n_155));
   AOI21_X1 i_220 (.A(n_163), .B1(n_159), .B2(n_158), .ZN(n_156));
   INV_X1 i_221 (.A(n_158), .ZN(n_157));
   NAND2_X1 i_222 (.A1(p_0[53]), .A2(adder[53]), .ZN(n_158));
   NAND2_X1 i_223 (.A1(p_0[52]), .A2(adder[52]), .ZN(n_159));
   NOR3_X1 i_224 (.A1(n_170), .A2(n_161), .A3(n_176), .ZN(n_160));
   OR2_X1 i_225 (.A1(n_163), .A2(n_162), .ZN(n_161));
   NOR2_X1 i_226 (.A1(p_0[52]), .A2(adder[52]), .ZN(n_162));
   NAND3_X1 i_227 (.A1(n_168), .A2(n_164), .A3(n_166), .ZN(n_163));
   INV_X1 i_228 (.A(n_165), .ZN(n_164));
   NOR2_X1 i_229 (.A1(p_0[54]), .A2(adder[54]), .ZN(n_165));
   INV_X1 i_230 (.A(n_167), .ZN(n_166));
   NOR2_X1 i_231 (.A1(p_0[53]), .A2(adder[53]), .ZN(n_167));
   INV_X1 i_232 (.A(n_169), .ZN(n_168));
   NOR2_X1 i_233 (.A1(p_0[55]), .A2(adder[55]), .ZN(n_169));
   OAI21_X1 i_234 (.A(n_171), .B1(p_0[56]), .B2(adder[56]), .ZN(n_170));
   NOR3_X1 i_235 (.A1(n_175), .A2(n_173), .A3(n_174), .ZN(n_171));
   NOR2_X1 i_236 (.A1(n_174), .A2(n_173), .ZN(n_172));
   NOR2_X1 i_237 (.A1(p_0[58]), .A2(adder[58]), .ZN(n_173));
   NOR2_X1 i_238 (.A1(p_0[57]), .A2(adder[57]), .ZN(n_174));
   NOR2_X1 i_239 (.A1(p_0[59]), .A2(adder[59]), .ZN(n_175));
   NOR4_X1 i_240 (.A1(n_180), .A2(n_177), .A3(n_181), .A4(n_184), .ZN(n_176));
   NOR2_X1 i_241 (.A1(n_189), .A2(n_179), .ZN(n_177));
   INV_X1 i_242 (.A(n_179), .ZN(n_178));
   NAND2_X1 i_243 (.A1(p_0[50]), .A2(adder[50]), .ZN(n_179));
   AND2_X1 i_244 (.A1(p_0[51]), .A2(adder[51]), .ZN(n_180));
   AOI21_X1 i_245 (.A(n_186), .B1(n_183), .B2(n_182), .ZN(n_181));
   NAND2_X1 i_246 (.A1(p_0[49]), .A2(adder[49]), .ZN(n_182));
   NAND2_X1 i_247 (.A1(p_0[48]), .A2(adder[48]), .ZN(n_183));
   NOR3_X1 i_248 (.A1(n_186), .A2(n_185), .A3(n_190), .ZN(n_184));
   NOR2_X1 i_249 (.A1(p_0[48]), .A2(adder[48]), .ZN(n_185));
   OR3_X1 i_250 (.A1(n_189), .A2(n_187), .A3(n_188), .ZN(n_186));
   NOR2_X1 i_251 (.A1(p_0[50]), .A2(adder[50]), .ZN(n_187));
   NOR2_X1 i_252 (.A1(p_0[49]), .A2(adder[49]), .ZN(n_188));
   NOR2_X1 i_253 (.A1(p_0[51]), .A2(adder[51]), .ZN(n_189));
   NOR3_X1 i_254 (.A1(n_212), .A2(n_191), .A3(n_219), .ZN(n_190));
   OAI221_X1 i_255 (.A(n_198), .B1(n_240), .B2(n_192), .C1(n_230), .C2(n_206), 
      .ZN(n_191));
   AOI221_X1 i_256 (.A(n_194), .B1(p_0[43]), .B2(adder[43]), .C1(n_238), 
      .C2(n_193), .ZN(n_192));
   AND2_X1 i_257 (.A1(p_0[42]), .A2(adder[42]), .ZN(n_193));
   AOI21_X1 i_258 (.A(n_233), .B1(n_197), .B2(n_196), .ZN(n_194));
   INV_X1 i_259 (.A(n_196), .ZN(n_195));
   NAND2_X1 i_260 (.A1(p_0[41]), .A2(adder[41]), .ZN(n_196));
   NAND2_X1 i_261 (.A1(p_0[40]), .A2(adder[40]), .ZN(n_197));
   AOI21_X1 i_262 (.A(n_199), .B1(p_0[47]), .B2(adder[47]), .ZN(n_198));
   OAI21_X1 i_263 (.A(n_202), .B1(n_245), .B2(n_201), .ZN(n_199));
   INV_X1 i_264 (.A(n_201), .ZN(n_200));
   NAND2_X1 i_265 (.A1(p_0[46]), .A2(adder[46]), .ZN(n_201));
   OAI21_X1 i_266 (.A(n_241), .B1(n_204), .B2(n_203), .ZN(n_202));
   AND2_X1 i_267 (.A1(p_0[45]), .A2(adder[45]), .ZN(n_203));
   INV_X1 i_268 (.A(n_205), .ZN(n_204));
   NAND2_X1 i_269 (.A1(p_0[44]), .A2(adder[44]), .ZN(n_205));
   AOI221_X1 i_270 (.A(n_208), .B1(p_0[39]), .B2(adder[39]), .C1(n_252), 
      .C2(n_207), .ZN(n_206));
   AND2_X1 i_271 (.A1(p_0[38]), .A2(adder[38]), .ZN(n_207));
   AOI21_X1 i_272 (.A(n_247), .B1(n_211), .B2(n_210), .ZN(n_208));
   INV_X1 i_273 (.A(n_210), .ZN(n_209));
   NAND2_X1 i_274 (.A1(p_0[37]), .A2(adder[37]), .ZN(n_210));
   NAND2_X1 i_275 (.A1(p_0[36]), .A2(adder[36]), .ZN(n_211));
   NOR2_X1 i_276 (.A1(n_229), .A2(n_213), .ZN(n_212));
   AOI221_X1 i_277 (.A(n_215), .B1(p_0[35]), .B2(adder[35]), .C1(n_227), 
      .C2(n_214), .ZN(n_213));
   AND2_X1 i_278 (.A1(p_0[34]), .A2(adder[34]), .ZN(n_214));
   AOI21_X1 i_279 (.A(n_222), .B1(n_218), .B2(n_217), .ZN(n_215));
   INV_X1 i_280 (.A(n_217), .ZN(n_216));
   NAND2_X1 i_281 (.A1(p_0[33]), .A2(adder[33]), .ZN(n_217));
   NAND2_X1 i_282 (.A1(p_0[32]), .A2(adder[32]), .ZN(n_218));
   NOR3_X1 i_283 (.A1(n_229), .A2(n_220), .A3(n_255), .ZN(n_219));
   OR2_X1 i_284 (.A1(n_222), .A2(n_221), .ZN(n_220));
   NOR2_X1 i_285 (.A1(p_0[32]), .A2(adder[32]), .ZN(n_221));
   NAND3_X1 i_286 (.A1(n_227), .A2(n_223), .A3(n_225), .ZN(n_222));
   INV_X1 i_287 (.A(n_224), .ZN(n_223));
   NOR2_X1 i_288 (.A1(p_0[34]), .A2(adder[34]), .ZN(n_224));
   INV_X1 i_289 (.A(n_226), .ZN(n_225));
   NOR2_X1 i_290 (.A1(p_0[33]), .A2(adder[33]), .ZN(n_226));
   INV_X1 i_291 (.A(n_228), .ZN(n_227));
   NOR2_X1 i_292 (.A1(p_0[35]), .A2(adder[35]), .ZN(n_228));
   OR2_X1 i_293 (.A1(n_246), .A2(n_230), .ZN(n_229));
   OR2_X1 i_294 (.A1(n_240), .A2(n_231), .ZN(n_230));
   OR2_X1 i_295 (.A1(n_233), .A2(n_232), .ZN(n_231));
   NOR2_X1 i_296 (.A1(p_0[40]), .A2(adder[40]), .ZN(n_232));
   NAND3_X1 i_297 (.A1(n_238), .A2(n_234), .A3(n_236), .ZN(n_233));
   INV_X1 i_298 (.A(n_235), .ZN(n_234));
   NOR2_X1 i_299 (.A1(p_0[42]), .A2(adder[42]), .ZN(n_235));
   INV_X1 i_300 (.A(n_237), .ZN(n_236));
   NOR2_X1 i_301 (.A1(p_0[41]), .A2(adder[41]), .ZN(n_237));
   INV_X1 i_302 (.A(n_239), .ZN(n_238));
   NOR2_X1 i_303 (.A1(p_0[43]), .A2(adder[43]), .ZN(n_239));
   OAI21_X1 i_304 (.A(n_241), .B1(p_0[44]), .B2(adder[44]), .ZN(n_240));
   NOR3_X1 i_305 (.A1(n_245), .A2(n_243), .A3(n_244), .ZN(n_241));
   NOR2_X1 i_306 (.A1(n_244), .A2(n_243), .ZN(n_242));
   NOR2_X1 i_307 (.A1(p_0[46]), .A2(adder[46]), .ZN(n_243));
   NOR2_X1 i_308 (.A1(p_0[45]), .A2(adder[45]), .ZN(n_244));
   NOR2_X1 i_309 (.A1(p_0[47]), .A2(adder[47]), .ZN(n_245));
   OR2_X1 i_310 (.A1(n_254), .A2(n_247), .ZN(n_246));
   NAND3_X1 i_311 (.A1(n_252), .A2(n_248), .A3(n_250), .ZN(n_247));
   INV_X1 i_312 (.A(n_249), .ZN(n_248));
   NOR2_X1 i_313 (.A1(p_0[38]), .A2(adder[38]), .ZN(n_249));
   INV_X1 i_314 (.A(n_251), .ZN(n_250));
   NOR2_X1 i_315 (.A1(p_0[37]), .A2(adder[37]), .ZN(n_251));
   INV_X1 i_316 (.A(n_253), .ZN(n_252));
   NOR2_X1 i_317 (.A1(p_0[39]), .A2(adder[39]), .ZN(n_253));
   NOR2_X1 i_318 (.A1(p_0[36]), .A2(adder[36]), .ZN(n_254));
   NOR3_X1 i_319 (.A1(n_263), .A2(n_256), .A3(n_281), .ZN(n_255));
   OAI222_X1 i_320 (.A1(n_291), .A2(n_275), .B1(n_292), .B2(n_257), .C1(n_302), 
      .C2(n_269), .ZN(n_256));
   AOI221_X1 i_321 (.A(n_259), .B1(p_0[23]), .B2(adder[23]), .C1(n_317), 
      .C2(n_258), .ZN(n_257));
   AND2_X1 i_322 (.A1(p_0[22]), .A2(adder[22]), .ZN(n_258));
   AOI21_X1 i_323 (.A(n_312), .B1(n_262), .B2(n_261), .ZN(n_259));
   INV_X1 i_324 (.A(n_261), .ZN(n_260));
   NAND2_X1 i_325 (.A1(p_0[21]), .A2(adder[21]), .ZN(n_261));
   NAND2_X1 i_326 (.A1(p_0[20]), .A2(adder[20]), .ZN(n_262));
   OAI222_X1 i_327 (.A1(n_304), .A2(n_266), .B1(n_310), .B2(n_265), .C1(n_377), 
      .C2(n_374), .ZN(n_263));
   INV_X1 i_328 (.A(n_265), .ZN(n_264));
   NAND2_X1 i_329 (.A1(p_0[30]), .A2(adder[30]), .ZN(n_265));
   AOI21_X1 i_330 (.A(n_267), .B1(p_0[28]), .B2(adder[28]), .ZN(n_266));
   AND2_X1 i_331 (.A1(p_0[29]), .A2(adder[29]), .ZN(n_267));
   NAND2_X1 i_332 (.A1(p_0[28]), .A2(adder[28]), .ZN(n_268));
   AOI221_X1 i_333 (.A(n_271), .B1(p_0[27]), .B2(adder[27]), .C1(n_300), 
      .C2(n_270), .ZN(n_269));
   AND2_X1 i_334 (.A1(p_0[26]), .A2(adder[26]), .ZN(n_270));
   AOI21_X1 i_335 (.A(n_295), .B1(n_274), .B2(n_273), .ZN(n_271));
   INV_X1 i_336 (.A(n_273), .ZN(n_272));
   NAND2_X1 i_337 (.A1(p_0[25]), .A2(adder[25]), .ZN(n_273));
   NAND2_X1 i_338 (.A1(p_0[24]), .A2(adder[24]), .ZN(n_274));
   AOI221_X1 i_339 (.A(n_277), .B1(p_0[19]), .B2(adder[19]), .C1(n_289), 
      .C2(n_276), .ZN(n_275));
   AND2_X1 i_340 (.A1(p_0[18]), .A2(adder[18]), .ZN(n_276));
   AOI21_X1 i_341 (.A(n_284), .B1(n_280), .B2(n_279), .ZN(n_277));
   INV_X1 i_342 (.A(n_279), .ZN(n_278));
   NAND2_X1 i_343 (.A1(p_0[17]), .A2(adder[17]), .ZN(n_279));
   NAND2_X1 i_344 (.A1(p_0[16]), .A2(adder[16]), .ZN(n_280));
   NOR3_X1 i_345 (.A1(n_291), .A2(n_282), .A3(n_320), .ZN(n_281));
   OR2_X1 i_346 (.A1(n_284), .A2(n_283), .ZN(n_282));
   NOR2_X1 i_347 (.A1(p_0[16]), .A2(adder[16]), .ZN(n_283));
   NAND3_X1 i_348 (.A1(n_289), .A2(n_285), .A3(n_287), .ZN(n_284));
   INV_X1 i_349 (.A(n_286), .ZN(n_285));
   NOR2_X1 i_350 (.A1(p_0[18]), .A2(adder[18]), .ZN(n_286));
   INV_X1 i_351 (.A(n_288), .ZN(n_287));
   NOR2_X1 i_352 (.A1(p_0[17]), .A2(adder[17]), .ZN(n_288));
   INV_X1 i_353 (.A(n_290), .ZN(n_289));
   NOR2_X1 i_354 (.A1(p_0[19]), .A2(adder[19]), .ZN(n_290));
   OR2_X1 i_355 (.A1(n_311), .A2(n_292), .ZN(n_291));
   OR2_X1 i_356 (.A1(n_302), .A2(n_293), .ZN(n_292));
   OR2_X1 i_357 (.A1(n_295), .A2(n_294), .ZN(n_293));
   NOR2_X1 i_358 (.A1(p_0[24]), .A2(adder[24]), .ZN(n_294));
   NAND3_X1 i_359 (.A1(n_300), .A2(n_296), .A3(n_298), .ZN(n_295));
   INV_X1 i_360 (.A(n_297), .ZN(n_296));
   NOR2_X1 i_361 (.A1(p_0[26]), .A2(adder[26]), .ZN(n_297));
   INV_X1 i_362 (.A(n_299), .ZN(n_298));
   NOR2_X1 i_363 (.A1(p_0[25]), .A2(adder[25]), .ZN(n_299));
   INV_X1 i_364 (.A(n_301), .ZN(n_300));
   NOR2_X1 i_365 (.A1(p_0[27]), .A2(adder[27]), .ZN(n_301));
   OR2_X1 i_366 (.A1(n_304), .A2(n_303), .ZN(n_302));
   NOR2_X1 i_367 (.A1(p_0[28]), .A2(adder[28]), .ZN(n_303));
   NAND3_X1 i_368 (.A1(n_309), .A2(n_305), .A3(n_307), .ZN(n_304));
   INV_X1 i_369 (.A(n_306), .ZN(n_305));
   NOR2_X1 i_370 (.A1(p_0[30]), .A2(adder[30]), .ZN(n_306));
   INV_X1 i_371 (.A(n_308), .ZN(n_307));
   NOR2_X1 i_372 (.A1(p_0[29]), .A2(adder[29]), .ZN(n_308));
   INV_X1 i_373 (.A(n_310), .ZN(n_309));
   NOR2_X1 i_374 (.A1(p_0[31]), .A2(adder[31]), .ZN(n_310));
   OR2_X1 i_375 (.A1(n_319), .A2(n_312), .ZN(n_311));
   NAND3_X1 i_376 (.A1(n_317), .A2(n_313), .A3(n_315), .ZN(n_312));
   INV_X1 i_377 (.A(n_314), .ZN(n_313));
   NOR2_X1 i_378 (.A1(p_0[22]), .A2(adder[22]), .ZN(n_314));
   INV_X1 i_379 (.A(n_316), .ZN(n_315));
   NOR2_X1 i_380 (.A1(p_0[21]), .A2(adder[21]), .ZN(n_316));
   INV_X1 i_381 (.A(n_318), .ZN(n_317));
   NOR2_X1 i_382 (.A1(p_0[23]), .A2(adder[23]), .ZN(n_318));
   NOR2_X1 i_383 (.A1(p_0[20]), .A2(adder[20]), .ZN(n_319));
   NOR4_X1 i_384 (.A1(n_324), .A2(n_321), .A3(n_325), .A4(n_328), .ZN(n_320));
   NOR2_X1 i_385 (.A1(n_333), .A2(n_323), .ZN(n_321));
   INV_X1 i_386 (.A(n_323), .ZN(n_322));
   NAND2_X1 i_387 (.A1(p_0[14]), .A2(adder[14]), .ZN(n_323));
   AND2_X1 i_388 (.A1(p_0[15]), .A2(adder[15]), .ZN(n_324));
   AOI21_X1 i_389 (.A(n_330), .B1(n_327), .B2(n_326), .ZN(n_325));
   NAND2_X1 i_390 (.A1(p_0[13]), .A2(adder[13]), .ZN(n_326));
   NAND2_X1 i_391 (.A1(p_0[12]), .A2(adder[12]), .ZN(n_327));
   NOR3_X1 i_392 (.A1(n_330), .A2(n_329), .A3(n_334), .ZN(n_328));
   NOR2_X1 i_393 (.A1(p_0[12]), .A2(adder[12]), .ZN(n_329));
   OR3_X1 i_394 (.A1(n_333), .A2(n_331), .A3(n_332), .ZN(n_330));
   NOR2_X1 i_395 (.A1(p_0[14]), .A2(adder[14]), .ZN(n_331));
   NOR2_X1 i_396 (.A1(p_0[13]), .A2(adder[13]), .ZN(n_332));
   NOR2_X1 i_397 (.A1(p_0[15]), .A2(adder[15]), .ZN(n_333));
   NOR4_X1 i_398 (.A1(n_338), .A2(n_335), .A3(n_339), .A4(n_342), .ZN(n_334));
   NOR2_X1 i_399 (.A1(n_347), .A2(n_337), .ZN(n_335));
   INV_X1 i_400 (.A(n_337), .ZN(n_336));
   NAND2_X1 i_401 (.A1(p_0[10]), .A2(adder[10]), .ZN(n_337));
   AND2_X1 i_402 (.A1(p_0[11]), .A2(adder[11]), .ZN(n_338));
   AOI21_X1 i_403 (.A(n_344), .B1(n_341), .B2(n_340), .ZN(n_339));
   NAND2_X1 i_404 (.A1(p_0[9]), .A2(adder[9]), .ZN(n_340));
   NAND2_X1 i_405 (.A1(p_0[8]), .A2(adder[8]), .ZN(n_341));
   NOR3_X1 i_406 (.A1(n_344), .A2(n_343), .A3(n_348), .ZN(n_342));
   NOR2_X1 i_407 (.A1(p_0[8]), .A2(adder[8]), .ZN(n_343));
   OR3_X1 i_408 (.A1(n_347), .A2(n_345), .A3(n_346), .ZN(n_344));
   NOR2_X1 i_409 (.A1(p_0[10]), .A2(adder[10]), .ZN(n_345));
   NOR2_X1 i_410 (.A1(p_0[9]), .A2(adder[9]), .ZN(n_346));
   NOR2_X1 i_411 (.A1(p_0[11]), .A2(adder[11]), .ZN(n_347));
   NOR4_X1 i_412 (.A1(n_352), .A2(n_349), .A3(n_353), .A4(n_356), .ZN(n_348));
   NOR2_X1 i_413 (.A1(n_361), .A2(n_351), .ZN(n_349));
   INV_X1 i_414 (.A(n_351), .ZN(n_350));
   NAND2_X1 i_415 (.A1(p_0[6]), .A2(adder[6]), .ZN(n_351));
   AND2_X1 i_416 (.A1(p_0[7]), .A2(adder[7]), .ZN(n_352));
   AOI21_X1 i_417 (.A(n_358), .B1(n_355), .B2(n_354), .ZN(n_353));
   NAND2_X1 i_418 (.A1(p_0[5]), .A2(adder[5]), .ZN(n_354));
   NAND2_X1 i_419 (.A1(p_0[4]), .A2(adder[4]), .ZN(n_355));
   NOR3_X1 i_420 (.A1(n_358), .A2(n_357), .A3(n_362), .ZN(n_356));
   NOR2_X1 i_421 (.A1(p_0[4]), .A2(adder[4]), .ZN(n_357));
   OR3_X1 i_422 (.A1(n_361), .A2(n_359), .A3(n_360), .ZN(n_358));
   NOR2_X1 i_423 (.A1(p_0[6]), .A2(adder[6]), .ZN(n_359));
   NOR2_X1 i_424 (.A1(p_0[5]), .A2(adder[5]), .ZN(n_360));
   NOR2_X1 i_425 (.A1(p_0[7]), .A2(adder[7]), .ZN(n_361));
   NAND2_X1 i_426 (.A1(n_371), .A2(n_363), .ZN(n_362));
   OAI21_X1 i_427 (.A(n_364), .B1(n_376), .B2(n_373), .ZN(n_363));
   OAI22_X1 i_428 (.A1(p_0[2]), .A2(adder[2]), .B1(n_369), .B2(n_365), .ZN(n_364));
   AOI21_X1 i_429 (.A(n_368), .B1(n_367), .B2(n_366), .ZN(n_365));
   NAND2_X1 i_430 (.A1(p_0[1]), .A2(adder[1]), .ZN(n_366));
   NAND2_X1 i_431 (.A1(p_0[0]), .A2(adder[0]), .ZN(n_367));
   NOR2_X1 i_432 (.A1(p_0[1]), .A2(adder[1]), .ZN(n_368));
   INV_X1 i_433 (.A(n_370), .ZN(n_369));
   NAND2_X1 i_434 (.A1(p_0[2]), .A2(adder[2]), .ZN(n_370));
   NAND2_X1 i_435 (.A1(n_376), .A2(n_373), .ZN(n_371));
   NOR2_X1 i_436 (.A1(p_0[60]), .A2(adder[60]), .ZN(n_372));
   INV_X1 i_437 (.A(adder[3]), .ZN(n_373));
   INV_X1 i_438 (.A(adder[31]), .ZN(n_374));
   INV_X1 i_439 (.A(adder[59]), .ZN(n_375));
   INV_X1 i_440 (.A(p_0[3]), .ZN(n_376));
   INV_X1 i_441 (.A(p_0[31]), .ZN(n_377));
   INV_X1 i_442 (.A(p_0[59]), .ZN(n_378));
endmodule

module Radix4_Booth_new(clk, rst, op1, op2, P);
   input clk;
   input rst;
   input [31:0]op1;
   input [31:0]op2;
   output [63:0]P;

   wire n_0_0;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_151;
   wire n_0_152;
   wire n_0_153;
   wire n_0_154;
   wire n_0_155;
   wire n_0_156;
   wire n_0_157;
   wire n_0_158;
   wire n_0_159;
   wire n_0_160;
   wire n_0_161;
   wire n_0_162;
   wire n_0_163;
   wire n_0_164;
   wire n_0_165;
   wire n_0_166;
   wire n_0_167;
   wire n_0_168;
   wire n_0_169;
   wire n_0_170;
   wire n_0_171;
   wire n_0_172;
   wire n_0_173;
   wire n_0_174;
   wire n_0_175;
   wire n_0_176;
   wire n_0_177;
   wire n_0_178;
   wire n_0_179;
   wire n_0_180;
   wire n_0_181;
   wire n_0_182;
   wire n_0_183;
   wire n_0_184;
   wire n_0_185;
   wire n_0_186;
   wire n_0_187;
   wire n_0_188;
   wire n_0_189;
   wire n_0_190;
   wire n_0_191;
   wire n_0_192;
   wire n_0_193;
   wire n_0_194;
   wire n_0_195;
   wire n_0_196;
   wire n_0_197;
   wire n_0_198;
   wire n_0_199;
   wire n_0_200;
   wire n_0_201;
   wire n_0_202;
   wire n_0_203;
   wire n_0_204;
   wire n_0_205;
   wire n_0_206;
   wire n_0_207;
   wire n_0_208;
   wire n_0_209;
   wire n_0_210;
   wire n_0_211;
   wire n_0_212;
   wire n_0_213;
   wire n_0_214;
   wire n_0_0_4;
   wire n_0_0_0;
   wire n_0_0_5;
   wire n_0_0_1;
   wire n_0_0_6;
   wire n_0_0_2;
   wire n_0_0_7;
   wire n_0_0_3;
   wire n_0_279;
   wire n_0_280;
   wire n_0_281;
   wire n_0_282;
   wire n_0_283;
   wire n_0_284;
   wire n_0_285;
   wire n_0_286;
   wire n_0_287;
   wire n_0_288;
   wire n_0_289;
   wire n_0_290;
   wire n_0_291;
   wire n_0_292;
   wire n_0_293;
   wire n_0_294;
   wire n_0_295;
   wire n_0_296;
   wire n_0_1;
   wire n_0_2;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_215;
   wire n_0_216;
   wire n_0_217;
   wire n_0_218;
   wire n_0_219;
   wire n_0_220;
   wire n_0_221;
   wire n_0_222;
   wire n_0_223;
   wire n_0_224;
   wire n_0_225;
   wire n_0_226;
   wire n_0_227;
   wire n_0_228;
   wire n_0_229;
   wire n_0_230;
   wire n_0_231;
   wire n_0_232;
   wire n_0_233;
   wire n_0_234;
   wire n_0_235;
   wire n_0_236;
   wire n_0_237;
   wire n_0_238;
   wire n_0_239;
   wire n_0_240;
   wire n_0_241;
   wire n_0_242;
   wire n_0_243;
   wire n_0_244;
   wire n_0_245;
   wire n_0_246;
   wire n_0_247;
   wire n_0_248;
   wire n_0_249;
   wire n_0_250;
   wire n_0_251;
   wire n_0_252;
   wire n_0_253;
   wire n_0_254;
   wire n_0_255;
   wire n_0_256;
   wire n_0_257;
   wire n_0_258;
   wire n_0_259;
   wire n_0_260;
   wire n_0_261;
   wire n_0_262;
   wire n_0_263;
   wire n_0_264;
   wire n_0_265;
   wire n_0_266;
   wire n_0_267;
   wire n_0_268;
   wire n_0_269;
   wire n_0_270;
   wire n_0_271;
   wire n_0_272;
   wire n_0_273;
   wire n_0_274;
   wire n_0_275;
   wire n_0_276;
   wire n_0_277;
   wire n_0_278;
   wire n_0_78;
   wire n_0_79;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_0_8;
   wire n_0_84;
   wire n_0_85;
   wire n_0_0_9;
   wire n_0_0_10;
   wire n_0_0_11;
   wire n_0_0_12;
   wire n_0_0_13;
   wire n_0_0_14;
   wire n_0_0_15;
   wire n_0_0_16;
   wire n_0_0_17;
   wire n_0_0_18;
   wire n_0_0_19;
   wire n_0_0_20;
   wire n_0_80;
   wire n_0_86;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_0_21;
   wire n_0_93;
   wire n_0_0_22;
   wire n_0_0_23;
   wire n_0_94;
   wire n_0_0_24;
   wire n_0_95;
   wire n_0_0_25;
   wire n_0_96;
   wire n_0_0_26;
   wire n_0_0_27;
   wire n_0_0_28;
   wire n_0_97;
   wire n_0_0_29;
   wire n_0_98;
   wire n_0_0_30;
   wire n_0_99;
   wire n_0_0_31;
   wire n_0_100;
   wire n_0_0_32;
   wire n_0_101;
   wire n_0_0_33;
   wire n_0_102;
   wire n_0_0_34;
   wire n_0_103;
   wire n_0_0_35;
   wire n_0_0_36;
   wire n_0_104;
   wire n_0_0_37;
   wire n_0_0_38;
   wire n_0_105;
   wire n_0_0_39;
   wire n_0_106;
   wire n_0_0_40;
   wire n_0_0_41;
   wire n_0_107;
   wire n_0_0_42;
   wire n_0_108;
   wire n_0_0_43;
   wire n_0_0_44;
   wire n_0_0_45;
   wire n_0_0_46;
   wire n_0_109;
   wire n_0_0_47;
   wire n_0_110;
   wire n_0_0_48;
   wire n_0_0_49;
   wire n_0_111;
   wire n_0_0_50;
   wire n_0_0_51;
   wire n_0_0_52;
   wire n_0_112;
   wire n_0_0_53;
   wire n_0_0_54;
   wire n_0_0_55;
   wire n_0_113;
   wire n_0_0_56;
   wire n_0_0_57;
   wire n_0_0_58;
   wire n_0_0_59;
   wire n_0_0_60;
   wire n_0_114;
   wire n_0_0_61;
   wire n_0_0_62;
   wire n_0_0_63;
   wire n_0_0_64;
   wire n_0_115;
   wire n_0_0_65;
   wire n_0_0_66;
   wire n_0_0_67;
   wire n_0_0_68;
   wire n_0_0_69;
   wire n_0_116;
   wire n_0_0_70;
   wire n_0_0_71;
   wire n_0_0_72;
   wire n_0_117;
   wire n_0_0_73;
   wire n_0_0_74;
   wire n_0_0_75;
   wire n_0_118;
   wire n_0_0_76;
   wire n_0_0_77;
   wire n_0_0_78;
   wire n_0_0_79;
   wire n_0_119;
   wire n_0_0_80;
   wire n_0_0_81;
   wire n_0_0_82;
   wire n_0_120;
   wire n_0_0_83;
   wire n_0_0_84;
   wire n_0_0_85;
   wire n_0_0_86;
   wire n_0_0_87;
   wire n_0_0_88;
   wire n_0_0_89;
   wire n_0_0_90;
   wire n_0_121;
   wire n_0_0_91;
   wire n_0_0_92;
   wire n_0_0_93;
   wire n_0_0_94;
   wire n_0_0_95;
   wire n_0_0_96;
   wire n_0_0_97;
   wire n_0_0_98;
   wire n_0_122;
   wire n_0_0_99;
   wire n_0_0_100;
   wire n_0_0_101;
   wire n_0_0_102;
   wire n_0_0_103;
   wire n_0_0_104;
   wire n_0_0_105;
   wire n_0_123;
   wire n_0_0_106;
   wire n_0_0_107;
   wire n_0_0_108;
   wire n_0_0_109;
   wire n_0_0_110;
   wire n_0_0_111;
   wire n_0_0_112;
   wire n_0_0_113;
   wire n_0_0_114;
   wire n_0_124;
   wire n_0_0_115;
   wire n_0_0_116;
   wire n_0_0_117;
   wire n_0_0_118;
   wire n_0_0_119;
   wire n_0_0_120;
   wire n_0_0_121;
   wire n_0_0_122;
   wire n_0_125;
   wire n_0_0_123;
   wire n_0_0_124;
   wire n_0_0_125;
   wire n_0_0_126;
   wire n_0_0_127;
   wire n_0_0_128;
   wire n_0_0_129;
   wire n_0_0_130;
   wire n_0_0_131;
   wire n_0_126;
   wire n_0_0_132;
   wire n_0_0_133;
   wire n_0_0_134;
   wire n_0_0_135;
   wire n_0_0_136;
   wire n_0_0_137;
   wire n_0_0_138;
   wire n_0_127;
   wire n_0_0_139;
   wire n_0_0_140;
   wire n_0_0_141;
   wire n_0_0_142;
   wire n_0_0_143;
   wire n_0_0_144;
   wire n_0_0_145;
   wire n_0_128;
   wire n_0_0_146;
   wire n_0_0_147;
   wire n_0_0_148;
   wire n_0_0_149;
   wire n_0_0_150;
   wire n_0_0_151;
   wire n_0_0_152;
   wire n_0_0_153;
   wire n_0_129;
   wire n_0_0_154;
   wire n_0_0_155;
   wire n_0_0_156;
   wire n_0_0_157;
   wire n_0_0_158;
   wire n_0_0_159;
   wire n_0_0_160;
   wire n_0_130;
   wire n_0_0_161;
   wire n_0_0_162;
   wire n_0_0_163;
   wire n_0_0_164;
   wire n_0_0_165;
   wire n_0_0_166;
   wire n_0_131;
   wire n_0_0_167;
   wire n_0_0_168;
   wire n_0_0_169;
   wire n_0_0_170;
   wire n_0_0_171;
   wire n_0_0_172;
   wire n_0_0_173;
   wire n_0_132;
   wire n_0_0_174;
   wire n_0_0_175;
   wire n_0_0_176;
   wire n_0_0_177;
   wire n_0_0_178;
   wire n_0_0_179;
   wire n_0_0_180;
   wire n_0_133;
   wire n_0_0_181;
   wire n_0_0_182;
   wire n_0_0_183;
   wire n_0_0_184;
   wire n_0_0_185;
   wire n_0_0_186;
   wire n_0_0_187;
   wire n_0_134;
   wire n_0_0_188;
   wire n_0_0_189;
   wire n_0_0_190;
   wire n_0_0_191;
   wire n_0_0_192;
   wire n_0_0_193;
   wire n_0_0_194;
   wire n_0_135;
   wire n_0_0_195;
   wire n_0_0_196;
   wire n_0_0_197;
   wire n_0_0_198;
   wire n_0_0_199;
   wire n_0_0_200;
   wire n_0_136;
   wire n_0_0_201;
   wire n_0_0_202;
   wire n_0_0_203;
   wire n_0_0_204;
   wire n_0_0_205;
   wire n_0_0_206;
   wire n_0_137;
   wire n_0_0_207;
   wire n_0_0_208;
   wire n_0_0_209;
   wire n_0_0_210;
   wire n_0_0_211;
   wire n_0_0_212;
   wire n_0_0_213;
   wire n_0_138;
   wire n_0_0_214;
   wire n_0_0_215;
   wire n_0_0_216;
   wire n_0_0_217;
   wire n_0_0_218;
   wire n_0_0_219;
   wire n_0_0_220;
   wire n_0_139;
   wire n_0_0_221;
   wire n_0_0_222;
   wire n_0_0_223;
   wire n_0_0_224;
   wire n_0_0_225;
   wire n_0_0_226;
   wire n_0_0_227;
   wire n_0_140;
   wire n_0_0_228;
   wire n_0_0_229;
   wire n_0_0_230;
   wire n_0_0_231;
   wire n_0_0_232;
   wire n_0_0_233;
   wire n_0_0_234;
   wire n_0_141;
   wire n_0_0_235;
   wire n_0_0_236;
   wire n_0_0_237;
   wire n_0_0_238;
   wire n_0_0_239;
   wire n_0_0_240;
   wire n_0_142;
   wire n_0_0_241;
   wire n_0_0_242;
   wire n_0_0_243;
   wire n_0_0_244;
   wire n_0_0_245;
   wire n_0_0_246;
   wire n_0_0_247;
   wire n_0_0_248;
   wire n_0_143;
   wire n_0_0_249;
   wire n_0_0_250;
   wire n_0_0_251;
   wire n_0_0_252;
   wire n_0_0_253;
   wire n_0_0_254;
   wire n_0_144;
   wire n_0_0_255;
   wire n_0_0_256;
   wire n_0_0_257;
   wire n_0_0_258;
   wire n_0_0_259;
   wire n_0_145;
   wire n_0_0_260;
   wire n_0_0_261;
   wire n_0_0_262;
   wire n_0_0_263;
   wire n_0_0_264;
   wire n_0_0_265;
   wire n_0_146;
   wire n_0_0_266;
   wire n_0_0_267;
   wire n_0_0_268;
   wire n_0_0_269;
   wire n_0_0_270;
   wire n_0_0_271;
   wire n_0_147;
   wire n_0_0_272;
   wire n_0_0_273;
   wire n_0_0_274;
   wire n_0_0_275;
   wire n_0_0_276;
   wire n_0_0_277;
   wire n_0_148;
   wire n_0_0_278;
   wire n_0_0_279;
   wire n_0_0_280;
   wire n_0_0_281;
   wire n_0_0_282;
   wire n_0_0_283;
   wire n_0_149;
   wire n_0_0_284;
   wire n_0_0_285;
   wire n_0_0_286;
   wire n_0_0_287;
   wire n_0_0_288;
   wire n_0_0_289;
   wire n_0_150;
   wire n_0_0_290;
   wire n_0_0_291;
   wire n_0_0_292;
   wire n_0_0_293;
   wire n_0_0_294;
   wire n_0_0_295;
   wire n_0_0_296;
   wire n_0_0_297;
   wire n_0_0_298;
   wire n_0_0_299;
   wire n_0_89;
   wire n_0_0_300;
   wire n_0_0_301;
   wire n_0_0_302;
   wire n_0_0_303;
   wire n_0_0_304;
   wire n_0_0_305;
   wire n_0_0_306;
   wire n_0_0_307;
   wire n_0_0_308;
   wire n_0_0_309;
   wire n_0_0_310;
   wire n_0_0_311;
   wire n_0_0_312;
   wire n_0_0_313;
   wire n_0_0_314;
   wire n_0_0_315;
   wire n_0_0_316;
   wire n_0_0_317;
   wire n_0_0_318;
   wire n_0_0_319;
   wire n_0_0_320;
   wire n_0_0_321;
   wire n_0_0_322;
   wire n_0_0_323;
   wire n_0_0_324;
   wire n_0_0_325;
   wire n_0_0_326;
   wire n_0_0_327;
   wire n_0_0_328;
   wire n_0_0_329;
   wire n_0_0_330;
   wire n_0_0_331;
   wire n_0_0_332;
   wire n_0_0_333;
   wire n_0_0_334;
   wire n_0_0_335;
   wire n_0_0_336;
   wire n_0_0_337;
   wire n_0_0_338;
   wire n_0_0_339;
   wire n_0_0_340;
   wire n_0_0_341;
   wire n_0_0_342;
   wire n_0_0_343;
   wire n_0_0_344;
   wire n_0_0_345;
   wire n_0_0_346;
   wire n_0_0_347;
   wire n_0_0_348;
   wire n_0_0_349;
   wire n_0_0_350;
   wire n_0_0_351;
   wire n_0_0_352;
   wire n_0_0_353;
   wire n_0_0_354;
   wire n_0_0_355;
   wire n_0_0_356;
   wire n_0_0_357;
   wire n_0_0_358;
   wire n_0_0_359;
   wire [63:0]adder;
   wire [5:0]n;
   wire n_0_87;
   wire [31:0]OP1_complement;
   wire q;
   wire n_0_88;

   CLKGATETST_X1 clk_gate_P_reg (.CK(clk), .E(n_0_86), .SE(1'b0), .GCK(n_0_0));
   DFF_X1 \P_reg[63]  (.D(n_0_77), .CK(n_0_0), .Q(P[63]), .QN());
   DFF_X1 \P_reg[62]  (.D(n_0_76), .CK(n_0_0), .Q(P[62]), .QN());
   DFF_X1 \P_reg[61]  (.D(n_0_75), .CK(n_0_0), .Q(P[61]), .QN());
   DFF_X1 \P_reg[60]  (.D(n_0_74), .CK(n_0_0), .Q(P[60]), .QN());
   DFF_X1 \P_reg[59]  (.D(n_0_73), .CK(n_0_0), .Q(P[59]), .QN());
   DFF_X1 \P_reg[58]  (.D(n_0_72), .CK(n_0_0), .Q(P[58]), .QN());
   DFF_X1 \P_reg[57]  (.D(n_0_71), .CK(n_0_0), .Q(P[57]), .QN());
   DFF_X1 \P_reg[56]  (.D(n_0_70), .CK(n_0_0), .Q(P[56]), .QN());
   DFF_X1 \P_reg[55]  (.D(n_0_69), .CK(n_0_0), .Q(P[55]), .QN());
   DFF_X1 \P_reg[54]  (.D(n_0_68), .CK(n_0_0), .Q(P[54]), .QN());
   DFF_X1 \P_reg[53]  (.D(n_0_67), .CK(n_0_0), .Q(P[53]), .QN());
   DFF_X1 \P_reg[52]  (.D(n_0_66), .CK(n_0_0), .Q(P[52]), .QN());
   DFF_X1 \P_reg[51]  (.D(n_0_65), .CK(n_0_0), .Q(P[51]), .QN());
   DFF_X1 \P_reg[50]  (.D(n_0_64), .CK(n_0_0), .Q(P[50]), .QN());
   DFF_X1 \P_reg[49]  (.D(n_0_63), .CK(n_0_0), .Q(P[49]), .QN());
   DFF_X1 \P_reg[48]  (.D(n_0_62), .CK(n_0_0), .Q(P[48]), .QN());
   DFF_X1 \P_reg[47]  (.D(n_0_61), .CK(n_0_0), .Q(P[47]), .QN());
   DFF_X1 \P_reg[46]  (.D(n_0_60), .CK(n_0_0), .Q(P[46]), .QN());
   DFF_X1 \P_reg[45]  (.D(n_0_59), .CK(n_0_0), .Q(P[45]), .QN());
   DFF_X1 \P_reg[44]  (.D(n_0_58), .CK(n_0_0), .Q(P[44]), .QN());
   DFF_X1 \P_reg[43]  (.D(n_0_57), .CK(n_0_0), .Q(P[43]), .QN());
   DFF_X1 \P_reg[42]  (.D(n_0_56), .CK(n_0_0), .Q(P[42]), .QN());
   DFF_X1 \P_reg[41]  (.D(n_0_55), .CK(n_0_0), .Q(P[41]), .QN());
   DFF_X1 \P_reg[40]  (.D(n_0_54), .CK(n_0_0), .Q(P[40]), .QN());
   DFF_X1 \P_reg[39]  (.D(n_0_53), .CK(n_0_0), .Q(P[39]), .QN());
   DFF_X1 \P_reg[38]  (.D(n_0_52), .CK(n_0_0), .Q(P[38]), .QN());
   DFF_X1 \P_reg[37]  (.D(n_0_51), .CK(n_0_0), .Q(P[37]), .QN());
   DFF_X1 \P_reg[36]  (.D(n_0_50), .CK(n_0_0), .Q(P[36]), .QN());
   DFF_X1 \P_reg[35]  (.D(n_0_49), .CK(n_0_0), .Q(P[35]), .QN());
   DFF_X1 \P_reg[34]  (.D(n_0_48), .CK(n_0_0), .Q(P[34]), .QN());
   DFF_X1 \P_reg[33]  (.D(n_0_47), .CK(n_0_0), .Q(P[33]), .QN());
   DFF_X1 \P_reg[32]  (.D(n_0_46), .CK(n_0_0), .Q(P[32]), .QN());
   DFF_X1 \P_reg[31]  (.D(n_0_45), .CK(n_0_0), .Q(P[31]), .QN());
   DFF_X1 \P_reg[30]  (.D(n_0_44), .CK(n_0_0), .Q(P[30]), .QN());
   DFF_X1 \P_reg[29]  (.D(n_0_43), .CK(n_0_0), .Q(P[29]), .QN());
   DFF_X1 \P_reg[28]  (.D(n_0_42), .CK(n_0_0), .Q(P[28]), .QN());
   DFF_X1 \P_reg[27]  (.D(n_0_41), .CK(n_0_0), .Q(P[27]), .QN());
   DFF_X1 \P_reg[26]  (.D(n_0_40), .CK(n_0_0), .Q(P[26]), .QN());
   DFF_X1 \P_reg[25]  (.D(n_0_39), .CK(n_0_0), .Q(P[25]), .QN());
   DFF_X1 \P_reg[24]  (.D(n_0_38), .CK(n_0_0), .Q(P[24]), .QN());
   DFF_X1 \P_reg[23]  (.D(n_0_37), .CK(n_0_0), .Q(P[23]), .QN());
   DFF_X1 \P_reg[22]  (.D(n_0_36), .CK(n_0_0), .Q(P[22]), .QN());
   DFF_X1 \P_reg[21]  (.D(n_0_35), .CK(n_0_0), .Q(P[21]), .QN());
   DFF_X1 \P_reg[20]  (.D(n_0_34), .CK(n_0_0), .Q(P[20]), .QN());
   DFF_X1 \P_reg[19]  (.D(n_0_2), .CK(n_0_0), .Q(P[19]), .QN());
   DFF_X1 \P_reg[18]  (.D(n_0_1), .CK(n_0_0), .Q(P[18]), .QN());
   DFF_X1 \P_reg[17]  (.D(n_0_296), .CK(n_0_0), .Q(P[17]), .QN());
   DFF_X1 \P_reg[16]  (.D(n_0_295), .CK(n_0_0), .Q(P[16]), .QN());
   DFF_X1 \P_reg[15]  (.D(n_0_294), .CK(n_0_0), .Q(P[15]), .QN());
   DFF_X1 \P_reg[14]  (.D(n_0_293), .CK(n_0_0), .Q(P[14]), .QN());
   DFF_X1 \P_reg[13]  (.D(n_0_292), .CK(n_0_0), .Q(P[13]), .QN());
   DFF_X1 \P_reg[12]  (.D(n_0_291), .CK(n_0_0), .Q(P[12]), .QN());
   DFF_X1 \P_reg[11]  (.D(n_0_290), .CK(n_0_0), .Q(P[11]), .QN());
   DFF_X1 \P_reg[10]  (.D(n_0_289), .CK(n_0_0), .Q(P[10]), .QN());
   DFF_X1 \P_reg[9]  (.D(n_0_288), .CK(n_0_0), .Q(P[9]), .QN());
   DFF_X1 \P_reg[8]  (.D(n_0_287), .CK(n_0_0), .Q(P[8]), .QN());
   DFF_X1 \P_reg[7]  (.D(n_0_286), .CK(n_0_0), .Q(P[7]), .QN());
   DFF_X1 \P_reg[6]  (.D(n_0_285), .CK(n_0_0), .Q(P[6]), .QN());
   DFF_X1 \P_reg[5]  (.D(n_0_284), .CK(n_0_0), .Q(P[5]), .QN());
   DFF_X1 \P_reg[4]  (.D(n_0_283), .CK(n_0_0), .Q(P[4]), .QN());
   DFF_X1 \P_reg[3]  (.D(n_0_282), .CK(n_0_0), .Q(P[3]), .QN());
   DFF_X1 \P_reg[2]  (.D(n_0_281), .CK(n_0_0), .Q(P[2]), .QN());
   DFF_X1 \P_reg[1]  (.D(n_0_280), .CK(n_0_0), .Q(P[1]), .QN());
   DFF_X1 \P_reg[0]  (.D(n_0_279), .CK(n_0_0), .Q(P[0]), .QN());
   datapath i_0_2 (.p_0({n_0_33, n_0_32, n_0_31, n_0_30, n_0_29, n_0_28, n_0_27, 
      n_0_26, n_0_25, n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, 
      n_0_17, n_0_16, n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, 
      n_0_8, n_0_7, n_0_6, n_0_5, n_0_4, n_0_3, uc_0}), .op1(op1));
   datapath__0_16 i_0_14 (.p_0({uc_1, uc_2, n_0_89, n_0_150, n_0_149, n_0_148, 
      n_0_147, n_0_146, n_0_145, n_0_144, n_0_143, n_0_142, n_0_141, n_0_140, 
      n_0_139, n_0_138, n_0_137, n_0_136, n_0_135, n_0_134, n_0_133, n_0_132, 
      n_0_131, n_0_130, n_0_129, n_0_128, n_0_127, n_0_126, n_0_125, n_0_124, 
      n_0_123, n_0_122, n_0_121, n_0_120, n_0_119, n_0_118, n_0_117, n_0_116, 
      n_0_115, n_0_114, n_0_113, n_0_112, n_0_111, n_0_110, n_0_109, n_0_108, 
      n_0_107, n_0_106, n_0_105, n_0_104, n_0_103, n_0_102, n_0_101, n_0_100, 
      n_0_99, n_0_98, n_0_97, n_0_96, n_0_95, n_0_94, n_0_93, n_0_92, n_0_91, 
      n_0_90}), .adder(adder), .p_1({n_0_214, n_0_213, n_0_212, n_0_211, n_0_210, 
      n_0_209, n_0_208, n_0_207, n_0_206, n_0_205, n_0_204, n_0_203, n_0_202, 
      n_0_201, n_0_200, n_0_199, n_0_198, n_0_197, n_0_196, n_0_195, n_0_194, 
      n_0_193, n_0_192, n_0_191, n_0_190, n_0_189, n_0_188, n_0_187, n_0_186, 
      n_0_185, n_0_184, n_0_183, n_0_182, n_0_181, n_0_180, n_0_179, n_0_178, 
      n_0_177, n_0_176, n_0_175, n_0_174, n_0_173, n_0_172, n_0_171, n_0_170, 
      n_0_169, n_0_168, n_0_167, n_0_166, n_0_165, n_0_164, n_0_163, n_0_162, 
      n_0_161, n_0_160, n_0_159, n_0_158, n_0_157, n_0_156, n_0_155, n_0_154, 
      n_0_153, n_0_152, n_0_151}));
   HA_X1 i_0_0_0 (.A(n[1]), .B(n[0]), .CO(n_0_0_0), .S(n_0_0_4));
   HA_X1 i_0_0_1 (.A(n[2]), .B(n_0_0_0), .CO(n_0_0_1), .S(n_0_0_5));
   HA_X1 i_0_0_2 (.A(n[3]), .B(n_0_0_1), .CO(n_0_0_2), .S(n_0_0_6));
   HA_X1 i_0_0_3 (.A(n[4]), .B(n_0_0_2), .CO(n_0_0_3), .S(n_0_0_7));
   AND2_X1 i_0_0_4 (.A1(n_0_0_354), .A2(adder[0]), .ZN(n_0_279));
   AND2_X1 i_0_0_5 (.A1(n_0_0_354), .A2(adder[1]), .ZN(n_0_280));
   AND2_X1 i_0_0_6 (.A1(n_0_0_354), .A2(adder[2]), .ZN(n_0_281));
   AND2_X1 i_0_0_7 (.A1(n_0_0_354), .A2(adder[3]), .ZN(n_0_282));
   AND2_X1 i_0_0_8 (.A1(n_0_0_354), .A2(adder[4]), .ZN(n_0_283));
   AND2_X1 i_0_0_9 (.A1(n_0_0_354), .A2(adder[5]), .ZN(n_0_284));
   AND2_X1 i_0_0_10 (.A1(n_0_0_354), .A2(adder[6]), .ZN(n_0_285));
   AND2_X1 i_0_0_11 (.A1(n_0_0_354), .A2(adder[7]), .ZN(n_0_286));
   AND2_X1 i_0_0_12 (.A1(n_0_0_354), .A2(adder[8]), .ZN(n_0_287));
   AND2_X1 i_0_0_13 (.A1(n_0_0_354), .A2(adder[9]), .ZN(n_0_288));
   AND2_X1 i_0_0_14 (.A1(n_0_0_354), .A2(adder[10]), .ZN(n_0_289));
   AND2_X1 i_0_0_15 (.A1(n_0_0_354), .A2(adder[11]), .ZN(n_0_290));
   AND2_X1 i_0_0_16 (.A1(n_0_0_354), .A2(adder[12]), .ZN(n_0_291));
   AND2_X1 i_0_0_17 (.A1(n_0_0_354), .A2(adder[13]), .ZN(n_0_292));
   AND2_X1 i_0_0_18 (.A1(n_0_0_354), .A2(adder[14]), .ZN(n_0_293));
   AND2_X1 i_0_0_19 (.A1(n_0_0_354), .A2(adder[15]), .ZN(n_0_294));
   AND2_X1 i_0_0_20 (.A1(n_0_0_354), .A2(adder[16]), .ZN(n_0_295));
   AND2_X1 i_0_0_21 (.A1(n_0_0_354), .A2(adder[17]), .ZN(n_0_296));
   AND2_X1 i_0_0_22 (.A1(n_0_0_354), .A2(adder[18]), .ZN(n_0_1));
   AND2_X1 i_0_0_23 (.A1(n_0_0_354), .A2(adder[19]), .ZN(n_0_2));
   AND2_X1 i_0_0_24 (.A1(n_0_0_354), .A2(adder[20]), .ZN(n_0_34));
   AND2_X1 i_0_0_25 (.A1(n_0_0_354), .A2(adder[21]), .ZN(n_0_35));
   AND2_X1 i_0_0_26 (.A1(n_0_0_354), .A2(adder[22]), .ZN(n_0_36));
   AND2_X1 i_0_0_27 (.A1(n_0_0_354), .A2(adder[23]), .ZN(n_0_37));
   AND2_X1 i_0_0_28 (.A1(n_0_0_354), .A2(adder[24]), .ZN(n_0_38));
   AND2_X1 i_0_0_29 (.A1(n_0_0_354), .A2(adder[25]), .ZN(n_0_39));
   AND2_X1 i_0_0_30 (.A1(n_0_0_354), .A2(adder[26]), .ZN(n_0_40));
   AND2_X1 i_0_0_31 (.A1(n_0_0_354), .A2(adder[27]), .ZN(n_0_41));
   AND2_X1 i_0_0_32 (.A1(n_0_0_354), .A2(adder[28]), .ZN(n_0_42));
   AND2_X1 i_0_0_33 (.A1(n_0_0_354), .A2(adder[29]), .ZN(n_0_43));
   AND2_X1 i_0_0_34 (.A1(n_0_0_354), .A2(adder[30]), .ZN(n_0_44));
   AND2_X1 i_0_0_35 (.A1(n_0_0_354), .A2(adder[31]), .ZN(n_0_45));
   AND2_X1 i_0_0_36 (.A1(n_0_0_354), .A2(adder[32]), .ZN(n_0_46));
   AND2_X1 i_0_0_37 (.A1(n_0_0_354), .A2(adder[33]), .ZN(n_0_47));
   AND2_X1 i_0_0_38 (.A1(n_0_0_354), .A2(adder[34]), .ZN(n_0_48));
   AND2_X1 i_0_0_39 (.A1(n_0_0_354), .A2(adder[35]), .ZN(n_0_49));
   AND2_X1 i_0_0_40 (.A1(n_0_0_354), .A2(adder[36]), .ZN(n_0_50));
   AND2_X1 i_0_0_41 (.A1(n_0_0_354), .A2(adder[37]), .ZN(n_0_51));
   AND2_X1 i_0_0_42 (.A1(n_0_0_354), .A2(adder[38]), .ZN(n_0_52));
   AND2_X1 i_0_0_43 (.A1(n_0_0_354), .A2(adder[39]), .ZN(n_0_53));
   AND2_X1 i_0_0_44 (.A1(n_0_0_354), .A2(adder[40]), .ZN(n_0_54));
   AND2_X1 i_0_0_45 (.A1(n_0_0_354), .A2(adder[41]), .ZN(n_0_55));
   AND2_X1 i_0_0_46 (.A1(n_0_0_354), .A2(adder[42]), .ZN(n_0_56));
   AND2_X1 i_0_0_47 (.A1(n_0_0_354), .A2(adder[43]), .ZN(n_0_57));
   AND2_X1 i_0_0_48 (.A1(n_0_0_354), .A2(adder[44]), .ZN(n_0_58));
   AND2_X1 i_0_0_49 (.A1(n_0_0_354), .A2(adder[45]), .ZN(n_0_59));
   AND2_X1 i_0_0_50 (.A1(n_0_0_354), .A2(adder[46]), .ZN(n_0_60));
   AND2_X1 i_0_0_51 (.A1(n_0_0_354), .A2(adder[47]), .ZN(n_0_61));
   AND2_X1 i_0_0_52 (.A1(n_0_0_354), .A2(adder[48]), .ZN(n_0_62));
   AND2_X1 i_0_0_53 (.A1(n_0_0_354), .A2(adder[49]), .ZN(n_0_63));
   AND2_X1 i_0_0_54 (.A1(n_0_0_354), .A2(adder[50]), .ZN(n_0_64));
   AND2_X1 i_0_0_55 (.A1(n_0_0_354), .A2(adder[51]), .ZN(n_0_65));
   AND2_X1 i_0_0_56 (.A1(n_0_0_354), .A2(adder[52]), .ZN(n_0_66));
   AND2_X1 i_0_0_57 (.A1(n_0_0_354), .A2(adder[53]), .ZN(n_0_67));
   AND2_X1 i_0_0_58 (.A1(n_0_0_354), .A2(adder[54]), .ZN(n_0_68));
   AND2_X1 i_0_0_59 (.A1(n_0_0_354), .A2(adder[55]), .ZN(n_0_69));
   AND2_X1 i_0_0_60 (.A1(n_0_0_354), .A2(adder[56]), .ZN(n_0_70));
   AND2_X1 i_0_0_61 (.A1(n_0_0_354), .A2(adder[57]), .ZN(n_0_71));
   AND2_X1 i_0_0_62 (.A1(n_0_0_354), .A2(adder[58]), .ZN(n_0_72));
   AND2_X1 i_0_0_63 (.A1(n_0_0_354), .A2(adder[59]), .ZN(n_0_73));
   AND2_X1 i_0_0_64 (.A1(n_0_0_354), .A2(adder[60]), .ZN(n_0_74));
   AND2_X1 i_0_0_65 (.A1(n_0_0_354), .A2(adder[61]), .ZN(n_0_75));
   AND2_X1 i_0_0_66 (.A1(n_0_0_354), .A2(adder[62]), .ZN(n_0_76));
   AND2_X1 i_0_0_67 (.A1(n_0_0_354), .A2(adder[63]), .ZN(n_0_77));
   AND2_X1 i_0_0_68 (.A1(n_0_0_354), .A2(n_0_151), .ZN(n_0_215));
   AND2_X1 i_0_0_69 (.A1(n_0_0_354), .A2(n_0_152), .ZN(n_0_216));
   AND2_X1 i_0_0_70 (.A1(n_0_0_354), .A2(n_0_153), .ZN(n_0_217));
   AND2_X1 i_0_0_71 (.A1(n_0_0_354), .A2(n_0_154), .ZN(n_0_218));
   AND2_X1 i_0_0_72 (.A1(n_0_0_354), .A2(n_0_155), .ZN(n_0_219));
   AND2_X1 i_0_0_73 (.A1(n_0_0_354), .A2(n_0_156), .ZN(n_0_220));
   AND2_X1 i_0_0_74 (.A1(n_0_0_354), .A2(n_0_157), .ZN(n_0_221));
   AND2_X1 i_0_0_75 (.A1(n_0_0_354), .A2(n_0_158), .ZN(n_0_222));
   AND2_X1 i_0_0_76 (.A1(n_0_0_354), .A2(n_0_159), .ZN(n_0_223));
   AND2_X1 i_0_0_77 (.A1(n_0_0_354), .A2(n_0_160), .ZN(n_0_224));
   AND2_X1 i_0_0_78 (.A1(n_0_0_354), .A2(n_0_161), .ZN(n_0_225));
   AND2_X1 i_0_0_79 (.A1(n_0_0_354), .A2(n_0_162), .ZN(n_0_226));
   AND2_X1 i_0_0_80 (.A1(n_0_0_354), .A2(n_0_163), .ZN(n_0_227));
   AND2_X1 i_0_0_81 (.A1(n_0_0_354), .A2(n_0_164), .ZN(n_0_228));
   AND2_X1 i_0_0_82 (.A1(n_0_0_354), .A2(n_0_165), .ZN(n_0_229));
   AND2_X1 i_0_0_83 (.A1(n_0_0_354), .A2(n_0_166), .ZN(n_0_230));
   AND2_X1 i_0_0_84 (.A1(n_0_0_354), .A2(n_0_167), .ZN(n_0_231));
   AND2_X1 i_0_0_85 (.A1(n_0_0_354), .A2(n_0_168), .ZN(n_0_232));
   AND2_X1 i_0_0_86 (.A1(n_0_0_354), .A2(n_0_169), .ZN(n_0_233));
   AND2_X1 i_0_0_87 (.A1(n_0_0_354), .A2(n_0_170), .ZN(n_0_234));
   AND2_X1 i_0_0_88 (.A1(n_0_0_354), .A2(n_0_171), .ZN(n_0_235));
   AND2_X1 i_0_0_89 (.A1(n_0_0_354), .A2(n_0_172), .ZN(n_0_236));
   AND2_X1 i_0_0_90 (.A1(n_0_0_354), .A2(n_0_173), .ZN(n_0_237));
   AND2_X1 i_0_0_91 (.A1(n_0_0_354), .A2(n_0_174), .ZN(n_0_238));
   AND2_X1 i_0_0_92 (.A1(n_0_0_354), .A2(n_0_175), .ZN(n_0_239));
   AND2_X1 i_0_0_93 (.A1(n_0_0_354), .A2(n_0_176), .ZN(n_0_240));
   AND2_X1 i_0_0_94 (.A1(n_0_0_354), .A2(n_0_177), .ZN(n_0_241));
   AND2_X1 i_0_0_95 (.A1(n_0_0_354), .A2(n_0_178), .ZN(n_0_242));
   AND2_X1 i_0_0_96 (.A1(n_0_0_354), .A2(n_0_179), .ZN(n_0_243));
   AND2_X1 i_0_0_97 (.A1(n_0_0_354), .A2(n_0_180), .ZN(n_0_244));
   AND2_X1 i_0_0_98 (.A1(n_0_0_354), .A2(n_0_181), .ZN(n_0_245));
   AND2_X1 i_0_0_99 (.A1(n_0_0_354), .A2(n_0_182), .ZN(n_0_246));
   AND2_X1 i_0_0_100 (.A1(n_0_0_354), .A2(n_0_183), .ZN(n_0_247));
   AND2_X1 i_0_0_101 (.A1(n_0_0_354), .A2(n_0_184), .ZN(n_0_248));
   AND2_X1 i_0_0_102 (.A1(n_0_0_354), .A2(n_0_185), .ZN(n_0_249));
   AND2_X1 i_0_0_103 (.A1(n_0_0_354), .A2(n_0_186), .ZN(n_0_250));
   AND2_X1 i_0_0_104 (.A1(n_0_0_354), .A2(n_0_187), .ZN(n_0_251));
   AND2_X1 i_0_0_105 (.A1(n_0_0_354), .A2(n_0_188), .ZN(n_0_252));
   AND2_X1 i_0_0_106 (.A1(n_0_0_354), .A2(n_0_189), .ZN(n_0_253));
   AND2_X1 i_0_0_107 (.A1(n_0_0_354), .A2(n_0_190), .ZN(n_0_254));
   AND2_X1 i_0_0_108 (.A1(n_0_0_354), .A2(n_0_191), .ZN(n_0_255));
   AND2_X1 i_0_0_109 (.A1(n_0_0_354), .A2(n_0_192), .ZN(n_0_256));
   AND2_X1 i_0_0_110 (.A1(n_0_0_354), .A2(n_0_193), .ZN(n_0_257));
   AND2_X1 i_0_0_111 (.A1(n_0_0_354), .A2(n_0_194), .ZN(n_0_258));
   AND2_X1 i_0_0_112 (.A1(n_0_0_354), .A2(n_0_195), .ZN(n_0_259));
   AND2_X1 i_0_0_113 (.A1(n_0_0_354), .A2(n_0_196), .ZN(n_0_260));
   AND2_X1 i_0_0_114 (.A1(n_0_0_354), .A2(n_0_197), .ZN(n_0_261));
   AND2_X1 i_0_0_115 (.A1(n_0_0_354), .A2(n_0_198), .ZN(n_0_262));
   AND2_X1 i_0_0_116 (.A1(n_0_0_354), .A2(n_0_199), .ZN(n_0_263));
   AND2_X1 i_0_0_117 (.A1(n_0_0_354), .A2(n_0_200), .ZN(n_0_264));
   AND2_X1 i_0_0_118 (.A1(n_0_0_354), .A2(n_0_201), .ZN(n_0_265));
   AND2_X1 i_0_0_119 (.A1(n_0_0_354), .A2(n_0_202), .ZN(n_0_266));
   AND2_X1 i_0_0_120 (.A1(n_0_0_354), .A2(n_0_203), .ZN(n_0_267));
   AND2_X1 i_0_0_121 (.A1(n_0_0_354), .A2(n_0_204), .ZN(n_0_268));
   AND2_X1 i_0_0_122 (.A1(n_0_0_354), .A2(n_0_205), .ZN(n_0_269));
   AND2_X1 i_0_0_123 (.A1(n_0_0_354), .A2(n_0_206), .ZN(n_0_270));
   AND2_X1 i_0_0_124 (.A1(n_0_0_354), .A2(n_0_207), .ZN(n_0_271));
   AND2_X1 i_0_0_125 (.A1(n_0_0_354), .A2(n_0_208), .ZN(n_0_272));
   AND2_X1 i_0_0_126 (.A1(n_0_0_354), .A2(n_0_209), .ZN(n_0_273));
   AND2_X1 i_0_0_127 (.A1(n_0_0_354), .A2(n_0_210), .ZN(n_0_274));
   AND2_X1 i_0_0_128 (.A1(n_0_0_354), .A2(n_0_211), .ZN(n_0_275));
   AND2_X1 i_0_0_129 (.A1(n_0_0_354), .A2(n_0_212), .ZN(n_0_276));
   AND2_X1 i_0_0_130 (.A1(n_0_0_354), .A2(n_0_213), .ZN(n_0_277));
   AND2_X1 i_0_0_131 (.A1(n_0_0_354), .A2(n_0_214), .ZN(n_0_278));
   NOR2_X1 i_0_0_132 (.A1(n[0]), .A2(rst), .ZN(n_0_78));
   NOR2_X1 i_0_0_133 (.A1(rst), .A2(n_0_0_353), .ZN(n_0_79));
   NOR2_X1 i_0_0_134 (.A1(rst), .A2(n_0_0_351), .ZN(n_0_81));
   AND2_X1 i_0_0_135 (.A1(n_0_0_354), .A2(n_0_0_7), .ZN(n_0_82));
   AOI211_X1 i_0_0_136 (.A(rst), .B(n_0_0_8), .C1(n[5]), .C2(n_0_0_3), .ZN(
      n_0_83));
   NOR2_X1 i_0_0_137 (.A1(n[5]), .A2(n_0_0_3), .ZN(n_0_0_8));
   OAI21_X1 i_0_0_138 (.A(n_0_0_354), .B1(n[5]), .B2(n[4]), .ZN(n_0_84));
   NAND2_X1 i_0_0_139 (.A1(n_0_0_15), .A2(n_0_0_9), .ZN(n_0_85));
   NAND3_X1 i_0_0_140 (.A1(n_0_0_354), .A2(n_0_0_352), .A3(n_0_0_10), .ZN(
      n_0_0_9));
   OAI33_X1 i_0_0_141 (.A1(n_0_0_351), .A2(n_0_0_13), .A3(n_0_0_14), .B1(
      n_0_0_12), .B2(n_0_0_11), .B3(n_0_0_6), .ZN(n_0_0_10));
   AOI221_X1 i_0_0_142 (.A(n_0_0_356), .B1(op2[3]), .B2(n_0_0_4), .C1(op2[31]), 
      .C2(n_0_0_353), .ZN(n_0_0_11));
   AOI221_X1 i_0_0_143 (.A(n[0]), .B1(op2[5]), .B2(n_0_0_4), .C1(op2[1]), 
      .C2(n_0_0_353), .ZN(n_0_0_12));
   AOI221_X1 i_0_0_144 (.A(n_0_0_4), .B1(n_0_0_356), .B2(op2[17]), .C1(n[0]), 
      .C2(op2[15]), .ZN(n_0_0_13));
   AOI221_X1 i_0_0_145 (.A(n_0_0_353), .B1(n_0_0_356), .B2(op2[21]), .C1(n[0]), 
      .C2(op2[19]), .ZN(n_0_0_14));
   NAND2_X1 i_0_0_146 (.A1(n_0_80), .A2(n_0_0_16), .ZN(n_0_0_15));
   OAI33_X1 i_0_0_147 (.A1(n_0_0_351), .A2(n_0_0_19), .A3(n_0_0_20), .B1(
      n_0_0_18), .B2(n_0_0_17), .B3(n_0_0_6), .ZN(n_0_0_16));
   AOI221_X1 i_0_0_148 (.A(n_0_0_356), .B1(op2[7]), .B2(n_0_0_353), .C1(op2[11]), 
      .C2(n_0_0_4), .ZN(n_0_0_17));
   AOI221_X1 i_0_0_149 (.A(n[0]), .B1(op2[9]), .B2(n_0_0_353), .C1(op2[13]), 
      .C2(n_0_0_4), .ZN(n_0_0_18));
   AOI221_X1 i_0_0_150 (.A(n_0_0_4), .B1(n_0_0_356), .B2(op2[25]), .C1(n[0]), 
      .C2(op2[23]), .ZN(n_0_0_19));
   AOI221_X1 i_0_0_151 (.A(n_0_0_353), .B1(n[0]), .B2(op2[27]), .C1(n_0_0_356), 
      .C2(op2[29]), .ZN(n_0_0_20));
   NOR2_X1 i_0_0_152 (.A1(rst), .A2(n_0_0_352), .ZN(n_0_80));
   OR3_X1 i_0_0_153 (.A1(n[5]), .A2(n[4]), .A3(rst), .ZN(n_0_86));
   AND2_X1 i_0_0_154 (.A1(n_0_0_89), .A2(n_0_0_23), .ZN(n_0_90));
   AND2_X1 i_0_0_155 (.A1(n_0_0_96), .A2(n_0_0_23), .ZN(n_0_91));
   INV_X1 i_0_0_156 (.A(n_0_0_21), .ZN(n_0_92));
   AOI22_X1 i_0_0_157 (.A1(n_0_0_103), .A2(n_0_0_23), .B1(n_0_0_338), .B2(
      n_0_0_89), .ZN(n_0_0_21));
   INV_X1 i_0_0_158 (.A(n_0_0_22), .ZN(n_0_93));
   AOI22_X1 i_0_0_159 (.A1(n_0_0_338), .A2(n_0_0_96), .B1(n_0_0_112), .B2(
      n_0_0_23), .ZN(n_0_0_22));
   NOR2_X1 i_0_0_160 (.A1(n[0]), .A2(n_0_0_315), .ZN(n_0_0_23));
   INV_X1 i_0_0_161 (.A(n_0_0_24), .ZN(n_0_94));
   AOI22_X1 i_0_0_162 (.A1(n_0_0_338), .A2(n_0_0_103), .B1(n_0_0_356), .B2(
      n_0_0_27), .ZN(n_0_0_24));
   OAI21_X1 i_0_0_163 (.A(n_0_0_25), .B1(n[0]), .B2(n_0_0_29), .ZN(n_0_95));
   NAND2_X1 i_0_0_164 (.A1(n_0_0_338), .A2(n_0_0_112), .ZN(n_0_0_25));
   OAI21_X1 i_0_0_165 (.A(n_0_0_26), .B1(n[0]), .B2(n_0_0_30), .ZN(n_0_96));
   NAND2_X1 i_0_0_166 (.A1(n[0]), .A2(n_0_0_27), .ZN(n_0_0_26));
   OAI21_X1 i_0_0_167 (.A(n_0_0_28), .B1(n_0_0_315), .B2(n_0_0_119), .ZN(
      n_0_0_27));
   NAND2_X1 i_0_0_168 (.A1(n_0_0_89), .A2(n_0_0_36), .ZN(n_0_0_28));
   OAI22_X1 i_0_0_169 (.A1(n[0]), .A2(n_0_0_31), .B1(n_0_0_356), .B2(n_0_0_29), 
      .ZN(n_0_97));
   AOI22_X1 i_0_0_170 (.A1(n_0_0_314), .A2(n_0_0_129), .B1(n_0_0_96), .B2(
      n_0_0_36), .ZN(n_0_0_29));
   OAI22_X1 i_0_0_171 (.A1(n[0]), .A2(n_0_0_32), .B1(n_0_0_356), .B2(n_0_0_30), 
      .ZN(n_0_98));
   AOI22_X1 i_0_0_172 (.A1(n_0_0_314), .A2(n_0_0_136), .B1(n_0_0_103), .B2(
      n_0_0_36), .ZN(n_0_0_30));
   OAI22_X1 i_0_0_173 (.A1(n[0]), .A2(n_0_0_33), .B1(n_0_0_356), .B2(n_0_0_31), 
      .ZN(n_0_99));
   AOI22_X1 i_0_0_174 (.A1(n_0_0_314), .A2(n_0_0_143), .B1(n_0_0_112), .B2(
      n_0_0_36), .ZN(n_0_0_31));
   OAI22_X1 i_0_0_175 (.A1(n[0]), .A2(n_0_0_34), .B1(n_0_0_356), .B2(n_0_0_32), 
      .ZN(n_0_100));
   AOI22_X1 i_0_0_176 (.A1(n_0_0_316), .A2(n_0_0_38), .B1(n_0_0_120), .B2(
      n_0_0_36), .ZN(n_0_0_32));
   OAI22_X1 i_0_0_177 (.A1(n[0]), .A2(n_0_0_35), .B1(n_0_0_356), .B2(n_0_0_33), 
      .ZN(n_0_101));
   AOI22_X1 i_0_0_178 (.A1(n_0_0_316), .A2(n_0_0_94), .B1(n_0_0_129), .B2(
      n_0_0_36), .ZN(n_0_0_33));
   OAI22_X1 i_0_0_179 (.A1(n[0]), .A2(n_0_0_37), .B1(n_0_0_356), .B2(n_0_0_34), 
      .ZN(n_0_102));
   AOI22_X1 i_0_0_180 (.A1(n_0_0_316), .A2(n_0_0_101), .B1(n_0_0_136), .B2(
      n_0_0_36), .ZN(n_0_0_34));
   OAI22_X1 i_0_0_181 (.A1(n[0]), .A2(n_0_0_39), .B1(n_0_0_356), .B2(n_0_0_35), 
      .ZN(n_0_103));
   AOI22_X1 i_0_0_182 (.A1(n_0_0_316), .A2(n_0_0_110), .B1(n_0_0_143), .B2(
      n_0_0_36), .ZN(n_0_0_35));
   NOR2_X1 i_0_0_183 (.A1(n_0_0_357), .A2(n_0_0_340), .ZN(n_0_0_36));
   OAI22_X1 i_0_0_184 (.A1(n[0]), .A2(n_0_0_41), .B1(n_0_0_356), .B2(n_0_0_37), 
      .ZN(n_0_104));
   AOI22_X1 i_0_0_185 (.A1(n_0_0_52), .A2(n_0_0_38), .B1(n_0_0_316), .B2(
      n_0_0_46), .ZN(n_0_0_37));
   AOI22_X1 i_0_0_186 (.A1(n_0_0_358), .A2(n_0_0_150), .B1(n[2]), .B2(n_0_0_90), 
      .ZN(n_0_0_38));
   OAI22_X1 i_0_0_187 (.A1(n[0]), .A2(n_0_0_42), .B1(n_0_0_356), .B2(n_0_0_39), 
      .ZN(n_0_105));
   AOI22_X1 i_0_0_188 (.A1(n_0_0_94), .A2(n_0_0_52), .B1(n_0_0_316), .B2(
      n_0_0_127), .ZN(n_0_0_39));
   OAI21_X1 i_0_0_189 (.A(n_0_0_40), .B1(n_0_0_356), .B2(n_0_0_41), .ZN(n_0_106));
   NAND2_X1 i_0_0_190 (.A1(n_0_0_356), .A2(n_0_0_44), .ZN(n_0_0_40));
   AOI22_X1 i_0_0_191 (.A1(n_0_0_101), .A2(n_0_0_52), .B1(n_0_0_316), .B2(
      n_0_0_134), .ZN(n_0_0_41));
   OAI22_X1 i_0_0_192 (.A1(n[0]), .A2(n_0_0_47), .B1(n_0_0_356), .B2(n_0_0_42), 
      .ZN(n_0_107));
   AOI22_X1 i_0_0_193 (.A1(n_0_0_110), .A2(n_0_0_52), .B1(n_0_0_316), .B2(
      n_0_0_141), .ZN(n_0_0_42));
   OAI21_X1 i_0_0_194 (.A(n_0_0_43), .B1(n[0]), .B2(n_0_0_49), .ZN(n_0_108));
   NAND2_X1 i_0_0_195 (.A1(n[0]), .A2(n_0_0_44), .ZN(n_0_0_43));
   OAI21_X1 i_0_0_196 (.A(n_0_0_45), .B1(n[1]), .B2(n_0_0_55), .ZN(n_0_0_44));
   NAND2_X1 i_0_0_197 (.A1(n_0_0_52), .A2(n_0_0_46), .ZN(n_0_0_45));
   AOI22_X1 i_0_0_198 (.A1(n[2]), .A2(n_0_0_119), .B1(n_0_0_358), .B2(n_0_0_177), 
      .ZN(n_0_0_46));
   OAI22_X1 i_0_0_199 (.A1(n[0]), .A2(n_0_0_51), .B1(n_0_0_356), .B2(n_0_0_47), 
      .ZN(n_0_109));
   AOI22_X1 i_0_0_200 (.A1(n_0_0_357), .A2(n_0_0_59), .B1(n_0_0_127), .B2(
      n_0_0_52), .ZN(n_0_0_47));
   OAI21_X1 i_0_0_201 (.A(n_0_0_48), .B1(n_0_0_356), .B2(n_0_0_49), .ZN(n_0_110));
   NAND2_X1 i_0_0_202 (.A1(n_0_0_356), .A2(n_0_0_54), .ZN(n_0_0_48));
   AOI22_X1 i_0_0_203 (.A1(n_0_0_357), .A2(n_0_0_63), .B1(n_0_0_134), .B2(
      n_0_0_52), .ZN(n_0_0_49));
   OAI21_X1 i_0_0_204 (.A(n_0_0_50), .B1(n_0_0_356), .B2(n_0_0_51), .ZN(n_0_111));
   NAND2_X1 i_0_0_205 (.A1(n_0_0_356), .A2(n_0_0_57), .ZN(n_0_0_50));
   AOI22_X1 i_0_0_206 (.A1(n_0_0_357), .A2(n_0_0_68), .B1(n_0_0_141), .B2(
      n_0_0_52), .ZN(n_0_0_51));
   NOR2_X1 i_0_0_207 (.A1(n[3]), .A2(n_0_0_357), .ZN(n_0_0_52));
   OAI21_X1 i_0_0_208 (.A(n_0_0_53), .B1(n[0]), .B2(n_0_0_62), .ZN(n_0_112));
   NAND2_X1 i_0_0_209 (.A1(n[0]), .A2(n_0_0_54), .ZN(n_0_0_53));
   AOI22_X1 i_0_0_210 (.A1(n_0_0_357), .A2(n_0_0_72), .B1(n[1]), .B2(n_0_0_55), 
      .ZN(n_0_0_54));
   AOI22_X1 i_0_0_211 (.A1(n_0_0_358), .A2(n_0_0_87), .B1(n_0_0_349), .B2(
      n_0_0_151), .ZN(n_0_0_55));
   INV_X1 i_0_0_212 (.A(n_0_0_56), .ZN(n_0_113));
   AOI22_X1 i_0_0_213 (.A1(n_0_0_356), .A2(n_0_0_66), .B1(n[0]), .B2(n_0_0_57), 
      .ZN(n_0_0_56));
   OAI21_X1 i_0_0_214 (.A(n_0_0_58), .B1(n[1]), .B2(n_0_0_75), .ZN(n_0_0_57));
   NAND2_X1 i_0_0_215 (.A1(n[1]), .A2(n_0_0_59), .ZN(n_0_0_58));
   OAI21_X1 i_0_0_216 (.A(n_0_0_60), .B1(n_0_0_340), .B2(n_0_0_210), .ZN(
      n_0_0_59));
   AOI22_X1 i_0_0_217 (.A1(n_0_0_349), .A2(n_0_0_158), .B1(n_0_0_342), .B2(
      n_0_0_96), .ZN(n_0_0_60));
   OAI21_X1 i_0_0_218 (.A(n_0_0_61), .B1(n_0_0_356), .B2(n_0_0_62), .ZN(n_0_114));
   NAND2_X1 i_0_0_219 (.A1(n_0_0_356), .A2(n_0_0_71), .ZN(n_0_0_61));
   AOI22_X1 i_0_0_220 (.A1(n[1]), .A2(n_0_0_63), .B1(n_0_0_357), .B2(n_0_0_78), 
      .ZN(n_0_0_62));
   OAI21_X1 i_0_0_221 (.A(n_0_0_64), .B1(n_0_0_340), .B2(n_0_0_217), .ZN(
      n_0_0_63));
   AOI22_X1 i_0_0_222 (.A1(n_0_0_349), .A2(n_0_0_164), .B1(n_0_0_342), .B2(
      n_0_0_103), .ZN(n_0_0_64));
   INV_X1 i_0_0_223 (.A(n_0_0_65), .ZN(n_0_115));
   AOI22_X1 i_0_0_224 (.A1(n_0_0_356), .A2(n_0_0_74), .B1(n[0]), .B2(n_0_0_66), 
      .ZN(n_0_0_65));
   OAI21_X1 i_0_0_225 (.A(n_0_0_67), .B1(n[1]), .B2(n_0_0_82), .ZN(n_0_0_66));
   NAND2_X1 i_0_0_226 (.A1(n[1]), .A2(n_0_0_68), .ZN(n_0_0_67));
   OAI21_X1 i_0_0_227 (.A(n_0_0_69), .B1(n_0_0_340), .B2(n_0_0_224), .ZN(
      n_0_0_68));
   AOI22_X1 i_0_0_228 (.A1(n_0_0_342), .A2(n_0_0_112), .B1(n_0_0_349), .B2(
      n_0_0_171), .ZN(n_0_0_69));
   OAI21_X1 i_0_0_229 (.A(n_0_0_70), .B1(n[0]), .B2(n_0_0_77), .ZN(n_0_116));
   NAND2_X1 i_0_0_230 (.A1(n[0]), .A2(n_0_0_71), .ZN(n_0_0_70));
   OAI22_X1 i_0_0_231 (.A1(n_0_0_357), .A2(n_0_0_72), .B1(n[1]), .B2(n_0_0_86), 
      .ZN(n_0_0_71));
   AOI22_X1 i_0_0_232 (.A1(n_0_0_358), .A2(n_0_0_118), .B1(n_0_0_349), .B2(
      n_0_0_178), .ZN(n_0_0_72));
   INV_X1 i_0_0_233 (.A(n_0_0_73), .ZN(n_0_117));
   AOI22_X1 i_0_0_234 (.A1(n[0]), .A2(n_0_0_74), .B1(n_0_0_356), .B2(n_0_0_81), 
      .ZN(n_0_0_73));
   AOI22_X1 i_0_0_235 (.A1(n_0_0_357), .A2(n_0_0_93), .B1(n[1]), .B2(n_0_0_75), 
      .ZN(n_0_0_74));
   AOI222_X1 i_0_0_236 (.A1(n_0_0_339), .A2(n_0_0_238), .B1(n_0_0_342), .B2(
      n_0_0_129), .C1(n_0_0_349), .C2(n_0_0_185), .ZN(n_0_0_75));
   OAI21_X1 i_0_0_237 (.A(n_0_0_76), .B1(n_0_0_356), .B2(n_0_0_77), .ZN(n_0_118));
   NAND2_X1 i_0_0_238 (.A1(n_0_0_356), .A2(n_0_0_84), .ZN(n_0_0_76));
   AOI22_X1 i_0_0_239 (.A1(n_0_0_357), .A2(n_0_0_100), .B1(n[1]), .B2(n_0_0_78), 
      .ZN(n_0_0_77));
   OAI21_X1 i_0_0_240 (.A(n_0_0_79), .B1(n_0_0_340), .B2(n_0_0_245), .ZN(
      n_0_0_78));
   AOI22_X1 i_0_0_241 (.A1(n_0_0_342), .A2(n_0_0_136), .B1(n_0_0_349), .B2(
      n_0_0_191), .ZN(n_0_0_79));
   INV_X1 i_0_0_242 (.A(n_0_0_80), .ZN(n_0_119));
   AOI22_X1 i_0_0_243 (.A1(n_0_0_356), .A2(n_0_0_92), .B1(n[0]), .B2(n_0_0_81), 
      .ZN(n_0_0_80));
   AOI22_X1 i_0_0_244 (.A1(n_0_0_357), .A2(n_0_0_109), .B1(n[1]), .B2(n_0_0_82), 
      .ZN(n_0_0_81));
   AOI222_X1 i_0_0_245 (.A1(n_0_0_339), .A2(n_0_0_252), .B1(n_0_0_342), .B2(
      n_0_0_143), .C1(n_0_0_349), .C2(n_0_0_198), .ZN(n_0_0_82));
   OAI21_X1 i_0_0_246 (.A(n_0_0_83), .B1(n[0]), .B2(n_0_0_99), .ZN(n_0_120));
   NAND2_X1 i_0_0_247 (.A1(n[0]), .A2(n_0_0_84), .ZN(n_0_0_83));
   OAI21_X1 i_0_0_248 (.A(n_0_0_85), .B1(n_0_0_357), .B2(n_0_0_86), .ZN(n_0_0_84));
   NAND2_X1 i_0_0_249 (.A1(n_0_0_357), .A2(n_0_0_116), .ZN(n_0_0_85));
   AOI22_X1 i_0_0_250 (.A1(n[2]), .A2(n_0_0_87), .B1(n_0_0_358), .B2(n_0_0_149), 
      .ZN(n_0_0_86));
   OAI21_X1 i_0_0_251 (.A(n_0_0_88), .B1(n_0_0_359), .B2(n_0_0_90), .ZN(n_0_0_87));
   NAND2_X1 i_0_0_252 (.A1(n_0_0_359), .A2(n_0_0_204), .ZN(n_0_0_88));
   INV_X1 i_0_0_253 (.A(n_0_0_90), .ZN(n_0_0_89));
   AOI22_X1 i_0_0_254 (.A1(OP1_complement[0]), .A2(n_0_0_304), .B1(op1[0]), 
      .B2(n_0_0_305), .ZN(n_0_0_90));
   INV_X1 i_0_0_255 (.A(n_0_0_91), .ZN(n_0_121));
   AOI22_X1 i_0_0_256 (.A1(n[0]), .A2(n_0_0_92), .B1(n_0_0_356), .B2(n_0_0_107), 
      .ZN(n_0_0_91));
   AOI22_X1 i_0_0_257 (.A1(n_0_0_357), .A2(n_0_0_126), .B1(n[1]), .B2(n_0_0_93), 
      .ZN(n_0_0_92));
   OAI222_X1 i_0_0_258 (.A1(n_0_0_340), .A2(n_0_0_263), .B1(n_0_0_350), .B2(
      n_0_0_211), .C1(n_0_0_359), .C2(n_0_0_94), .ZN(n_0_0_93));
   AOI21_X1 i_0_0_259 (.A(n_0_0_95), .B1(n_0_0_358), .B2(n_0_0_157), .ZN(
      n_0_0_94));
   NOR2_X1 i_0_0_260 (.A1(n_0_0_358), .A2(n_0_0_96), .ZN(n_0_0_95));
   NAND2_X1 i_0_0_261 (.A1(n_0_0_98), .A2(n_0_0_97), .ZN(n_0_0_96));
   AOI22_X1 i_0_0_262 (.A1(op1[1]), .A2(n_0_0_305), .B1(op1[0]), .B2(n_0_0_303), 
      .ZN(n_0_0_97));
   AOI22_X1 i_0_0_263 (.A1(OP1_complement[1]), .A2(n_0_0_304), .B1(
      OP1_complement[0]), .B2(n_0_0_302), .ZN(n_0_0_98));
   OAI22_X1 i_0_0_264 (.A1(n[0]), .A2(n_0_0_115), .B1(n_0_0_356), .B2(n_0_0_99), 
      .ZN(n_0_122));
   AOI22_X1 i_0_0_265 (.A1(n[1]), .A2(n_0_0_100), .B1(n_0_0_357), .B2(n_0_0_133), 
      .ZN(n_0_0_99));
   AOI222_X1 i_0_0_266 (.A1(n_0_0_339), .A2(n_0_0_268), .B1(n_0_0_349), .B2(
      n_0_0_217), .C1(n[3]), .C2(n_0_0_102), .ZN(n_0_0_100));
   INV_X1 i_0_0_267 (.A(n_0_0_102), .ZN(n_0_0_101));
   OAI22_X1 i_0_0_268 (.A1(n_0_0_358), .A2(n_0_0_103), .B1(n[2]), .B2(n_0_0_164), 
      .ZN(n_0_0_102));
   NAND2_X1 i_0_0_269 (.A1(n_0_0_105), .A2(n_0_0_104), .ZN(n_0_0_103));
   AOI22_X1 i_0_0_270 (.A1(op1[2]), .A2(n_0_0_305), .B1(op1[1]), .B2(n_0_0_303), 
      .ZN(n_0_0_104));
   AOI22_X1 i_0_0_271 (.A1(OP1_complement[2]), .A2(n_0_0_304), .B1(
      OP1_complement[1]), .B2(n_0_0_302), .ZN(n_0_0_105));
   INV_X1 i_0_0_272 (.A(n_0_0_106), .ZN(n_0_123));
   AOI22_X1 i_0_0_273 (.A1(n_0_0_356), .A2(n_0_0_124), .B1(n[0]), .B2(n_0_0_107), 
      .ZN(n_0_0_106));
   OAI21_X1 i_0_0_274 (.A(n_0_0_108), .B1(n_0_0_357), .B2(n_0_0_109), .ZN(
      n_0_0_107));
   NAND2_X1 i_0_0_275 (.A1(n_0_0_357), .A2(n_0_0_140), .ZN(n_0_0_108));
   OAI222_X1 i_0_0_276 (.A1(n_0_0_350), .A2(n_0_0_225), .B1(n_0_0_340), .B2(
      n_0_0_275), .C1(n_0_0_359), .C2(n_0_0_110), .ZN(n_0_0_109));
   AOI21_X1 i_0_0_277 (.A(n_0_0_111), .B1(n_0_0_358), .B2(n_0_0_170), .ZN(
      n_0_0_110));
   NOR2_X1 i_0_0_278 (.A1(n_0_0_358), .A2(n_0_0_112), .ZN(n_0_0_111));
   NAND2_X1 i_0_0_279 (.A1(n_0_0_114), .A2(n_0_0_113), .ZN(n_0_0_112));
   AOI22_X1 i_0_0_280 (.A1(op1[3]), .A2(n_0_0_305), .B1(op1[2]), .B2(n_0_0_303), 
      .ZN(n_0_0_113));
   AOI22_X1 i_0_0_281 (.A1(OP1_complement[3]), .A2(n_0_0_304), .B1(
      OP1_complement[2]), .B2(n_0_0_302), .ZN(n_0_0_114));
   OAI22_X1 i_0_0_282 (.A1(n_0_0_356), .A2(n_0_0_115), .B1(n[0]), .B2(n_0_0_132), 
      .ZN(n_0_124));
   AOI22_X1 i_0_0_283 (.A1(n[1]), .A2(n_0_0_116), .B1(n_0_0_357), .B2(n_0_0_147), 
      .ZN(n_0_0_115));
   AOI222_X1 i_0_0_284 (.A1(n_0_0_339), .A2(n_0_0_280), .B1(n_0_0_342), .B2(
      n_0_0_177), .C1(n[2]), .C2(n_0_0_117), .ZN(n_0_0_116));
   INV_X1 i_0_0_285 (.A(n_0_0_118), .ZN(n_0_0_117));
   AOI22_X1 i_0_0_286 (.A1(n_0_0_359), .A2(n_0_0_231), .B1(n[3]), .B2(n_0_0_119), 
      .ZN(n_0_0_118));
   INV_X1 i_0_0_287 (.A(n_0_0_120), .ZN(n_0_0_119));
   NAND2_X1 i_0_0_288 (.A1(n_0_0_122), .A2(n_0_0_121), .ZN(n_0_0_120));
   AOI22_X1 i_0_0_289 (.A1(op1[4]), .A2(n_0_0_305), .B1(OP1_complement[4]), 
      .B2(n_0_0_304), .ZN(n_0_0_121));
   AOI22_X1 i_0_0_290 (.A1(op1[3]), .A2(n_0_0_303), .B1(OP1_complement[3]), 
      .B2(n_0_0_302), .ZN(n_0_0_122));
   OAI21_X1 i_0_0_291 (.A(n_0_0_123), .B1(n[0]), .B2(n_0_0_139), .ZN(n_0_125));
   NAND2_X1 i_0_0_292 (.A1(n[0]), .A2(n_0_0_124), .ZN(n_0_0_123));
   OAI21_X1 i_0_0_293 (.A(n_0_0_125), .B1(n_0_0_357), .B2(n_0_0_126), .ZN(
      n_0_0_124));
   NAND2_X1 i_0_0_294 (.A1(n_0_0_357), .A2(n_0_0_155), .ZN(n_0_0_125));
   OAI222_X1 i_0_0_295 (.A1(n_0_0_340), .A2(n_0_0_287), .B1(n_0_0_350), .B2(
      n_0_0_238), .C1(n_0_0_359), .C2(n_0_0_127), .ZN(n_0_0_126));
   AOI21_X1 i_0_0_296 (.A(n_0_0_128), .B1(n_0_0_358), .B2(n_0_0_184), .ZN(
      n_0_0_127));
   NOR2_X1 i_0_0_297 (.A1(n_0_0_358), .A2(n_0_0_129), .ZN(n_0_0_128));
   NAND2_X1 i_0_0_298 (.A1(n_0_0_131), .A2(n_0_0_130), .ZN(n_0_0_129));
   AOI22_X1 i_0_0_299 (.A1(op1[5]), .A2(n_0_0_305), .B1(op1[4]), .B2(n_0_0_303), 
      .ZN(n_0_0_130));
   AOI22_X1 i_0_0_300 (.A1(OP1_complement[5]), .A2(n_0_0_304), .B1(
      OP1_complement[4]), .B2(n_0_0_302), .ZN(n_0_0_131));
   OAI22_X1 i_0_0_301 (.A1(n_0_0_356), .A2(n_0_0_132), .B1(n[0]), .B2(n_0_0_146), 
      .ZN(n_0_126));
   AOI22_X1 i_0_0_302 (.A1(n[1]), .A2(n_0_0_133), .B1(n_0_0_357), .B2(n_0_0_162), 
      .ZN(n_0_0_132));
   AOI222_X1 i_0_0_303 (.A1(n_0_0_339), .A2(n_0_0_292), .B1(n_0_0_349), .B2(
      n_0_0_245), .C1(n[3]), .C2(n_0_0_135), .ZN(n_0_0_133));
   INV_X1 i_0_0_304 (.A(n_0_0_135), .ZN(n_0_0_134));
   OAI22_X1 i_0_0_305 (.A1(n_0_0_358), .A2(n_0_0_136), .B1(n[2]), .B2(n_0_0_191), 
      .ZN(n_0_0_135));
   NAND2_X1 i_0_0_306 (.A1(n_0_0_138), .A2(n_0_0_137), .ZN(n_0_0_136));
   AOI22_X1 i_0_0_307 (.A1(op1[6]), .A2(n_0_0_305), .B1(OP1_complement[6]), 
      .B2(n_0_0_304), .ZN(n_0_0_137));
   AOI22_X1 i_0_0_308 (.A1(op1[5]), .A2(n_0_0_303), .B1(OP1_complement[5]), 
      .B2(n_0_0_302), .ZN(n_0_0_138));
   OAI22_X1 i_0_0_309 (.A1(n_0_0_356), .A2(n_0_0_139), .B1(n[0]), .B2(n_0_0_154), 
      .ZN(n_0_127));
   AOI22_X1 i_0_0_310 (.A1(n_0_0_357), .A2(n_0_0_168), .B1(n[1]), .B2(n_0_0_140), 
      .ZN(n_0_0_139));
   AOI221_X1 i_0_0_311 (.A(n_0_0_194), .B1(n_0_0_349), .B2(n_0_0_251), .C1(n[3]), 
      .C2(n_0_0_142), .ZN(n_0_0_140));
   INV_X1 i_0_0_312 (.A(n_0_0_142), .ZN(n_0_0_141));
   OAI22_X1 i_0_0_313 (.A1(n_0_0_358), .A2(n_0_0_143), .B1(n[2]), .B2(n_0_0_198), 
      .ZN(n_0_0_142));
   NAND2_X1 i_0_0_314 (.A1(n_0_0_145), .A2(n_0_0_144), .ZN(n_0_0_143));
   AOI22_X1 i_0_0_315 (.A1(op1[7]), .A2(n_0_0_305), .B1(OP1_complement[7]), 
      .B2(n_0_0_304), .ZN(n_0_0_144));
   AOI22_X1 i_0_0_316 (.A1(op1[6]), .A2(n_0_0_303), .B1(OP1_complement[6]), 
      .B2(n_0_0_302), .ZN(n_0_0_145));
   OAI22_X1 i_0_0_317 (.A1(n[0]), .A2(n_0_0_161), .B1(n_0_0_356), .B2(n_0_0_146), 
      .ZN(n_0_128));
   AOI22_X1 i_0_0_318 (.A1(n_0_0_357), .A2(n_0_0_175), .B1(n[1]), .B2(n_0_0_147), 
      .ZN(n_0_0_146));
   OAI21_X1 i_0_0_319 (.A(n_0_0_148), .B1(n_0_0_340), .B2(n_0_0_299), .ZN(
      n_0_0_147));
   AOI22_X1 i_0_0_320 (.A1(n[2]), .A2(n_0_0_149), .B1(n_0_0_342), .B2(n_0_0_204), 
      .ZN(n_0_0_148));
   AOI22_X1 i_0_0_321 (.A1(n_0_0_359), .A2(n_0_0_257), .B1(n[3]), .B2(n_0_0_150), 
      .ZN(n_0_0_149));
   INV_X1 i_0_0_322 (.A(n_0_0_151), .ZN(n_0_0_150));
   NAND2_X1 i_0_0_323 (.A1(n_0_0_153), .A2(n_0_0_152), .ZN(n_0_0_151));
   AOI22_X1 i_0_0_324 (.A1(op1[8]), .A2(n_0_0_305), .B1(op1[7]), .B2(n_0_0_303), 
      .ZN(n_0_0_152));
   AOI22_X1 i_0_0_325 (.A1(OP1_complement[8]), .A2(n_0_0_304), .B1(
      OP1_complement[7]), .B2(n_0_0_302), .ZN(n_0_0_153));
   OAI22_X1 i_0_0_326 (.A1(n[0]), .A2(n_0_0_167), .B1(n_0_0_356), .B2(n_0_0_154), 
      .ZN(n_0_129));
   AOI22_X1 i_0_0_327 (.A1(n_0_0_357), .A2(n_0_0_182), .B1(n[1]), .B2(n_0_0_155), 
      .ZN(n_0_0_154));
   AOI211_X1 i_0_0_328 (.A(n_0_0_194), .B(n_0_0_156), .C1(n_0_0_344), .C2(
      n_0_0_157), .ZN(n_0_0_155));
   OAI22_X1 i_0_0_329 (.A1(n_0_0_343), .A2(n_0_0_211), .B1(n_0_0_350), .B2(
      n_0_0_263), .ZN(n_0_0_156));
   INV_X1 i_0_0_330 (.A(n_0_0_158), .ZN(n_0_0_157));
   NAND2_X1 i_0_0_331 (.A1(n_0_0_160), .A2(n_0_0_159), .ZN(n_0_0_158));
   AOI22_X1 i_0_0_332 (.A1(op1[9]), .A2(n_0_0_305), .B1(op1[8]), .B2(n_0_0_303), 
      .ZN(n_0_0_159));
   AOI22_X1 i_0_0_333 (.A1(OP1_complement[9]), .A2(n_0_0_304), .B1(
      OP1_complement[8]), .B2(n_0_0_302), .ZN(n_0_0_160));
   OAI22_X1 i_0_0_334 (.A1(n[0]), .A2(n_0_0_174), .B1(n_0_0_356), .B2(n_0_0_161), 
      .ZN(n_0_130));
   AOI22_X1 i_0_0_335 (.A1(n_0_0_357), .A2(n_0_0_189), .B1(n[1]), .B2(n_0_0_162), 
      .ZN(n_0_0_161));
   AOI211_X1 i_0_0_336 (.A(n_0_0_194), .B(n_0_0_163), .C1(n_0_0_349), .C2(
      n_0_0_268), .ZN(n_0_0_162));
   OAI22_X1 i_0_0_337 (.A1(n_0_0_343), .A2(n_0_0_218), .B1(n_0_0_345), .B2(
      n_0_0_164), .ZN(n_0_0_163));
   NAND2_X1 i_0_0_338 (.A1(n_0_0_166), .A2(n_0_0_165), .ZN(n_0_0_164));
   AOI22_X1 i_0_0_339 (.A1(op1[10]), .A2(n_0_0_305), .B1(op1[9]), .B2(n_0_0_303), 
      .ZN(n_0_0_165));
   AOI22_X1 i_0_0_340 (.A1(OP1_complement[10]), .A2(n_0_0_304), .B1(
      OP1_complement[9]), .B2(n_0_0_302), .ZN(n_0_0_166));
   OAI22_X1 i_0_0_341 (.A1(n_0_0_356), .A2(n_0_0_167), .B1(n[0]), .B2(n_0_0_181), 
      .ZN(n_0_131));
   AOI22_X1 i_0_0_342 (.A1(n[1]), .A2(n_0_0_168), .B1(n_0_0_357), .B2(n_0_0_196), 
      .ZN(n_0_0_167));
   AOI211_X1 i_0_0_343 (.A(n_0_0_194), .B(n_0_0_169), .C1(n_0_0_344), .C2(
      n_0_0_170), .ZN(n_0_0_168));
   OAI22_X1 i_0_0_344 (.A1(n_0_0_350), .A2(n_0_0_275), .B1(n_0_0_343), .B2(
      n_0_0_225), .ZN(n_0_0_169));
   INV_X1 i_0_0_345 (.A(n_0_0_171), .ZN(n_0_0_170));
   NAND2_X1 i_0_0_346 (.A1(n_0_0_173), .A2(n_0_0_172), .ZN(n_0_0_171));
   AOI22_X1 i_0_0_347 (.A1(op1[11]), .A2(n_0_0_305), .B1(op1[10]), .B2(n_0_0_303), 
      .ZN(n_0_0_172));
   AOI22_X1 i_0_0_348 (.A1(OP1_complement[11]), .A2(n_0_0_304), .B1(
      OP1_complement[10]), .B2(n_0_0_302), .ZN(n_0_0_173));
   OAI22_X1 i_0_0_349 (.A1(n_0_0_356), .A2(n_0_0_174), .B1(n[0]), .B2(n_0_0_188), 
      .ZN(n_0_132));
   AOI22_X1 i_0_0_350 (.A1(n[1]), .A2(n_0_0_175), .B1(n_0_0_357), .B2(n_0_0_202), 
      .ZN(n_0_0_174));
   AOI211_X1 i_0_0_351 (.A(n_0_0_194), .B(n_0_0_176), .C1(n_0_0_349), .C2(
      n_0_0_280), .ZN(n_0_0_175));
   OAI22_X1 i_0_0_352 (.A1(n_0_0_343), .A2(n_0_0_232), .B1(n_0_0_345), .B2(
      n_0_0_178), .ZN(n_0_0_176));
   INV_X1 i_0_0_353 (.A(n_0_0_178), .ZN(n_0_0_177));
   NAND2_X1 i_0_0_354 (.A1(n_0_0_180), .A2(n_0_0_179), .ZN(n_0_0_178));
   AOI22_X1 i_0_0_355 (.A1(OP1_complement[12]), .A2(n_0_0_304), .B1(op1[11]), 
      .B2(n_0_0_303), .ZN(n_0_0_179));
   AOI22_X1 i_0_0_356 (.A1(op1[12]), .A2(n_0_0_305), .B1(OP1_complement[11]), 
      .B2(n_0_0_302), .ZN(n_0_0_180));
   OAI22_X1 i_0_0_357 (.A1(n_0_0_356), .A2(n_0_0_181), .B1(n[0]), .B2(n_0_0_195), 
      .ZN(n_0_133));
   AOI22_X1 i_0_0_358 (.A1(n[1]), .A2(n_0_0_182), .B1(n_0_0_357), .B2(n_0_0_208), 
      .ZN(n_0_0_181));
   AOI211_X1 i_0_0_359 (.A(n_0_0_194), .B(n_0_0_183), .C1(n_0_0_344), .C2(
      n_0_0_184), .ZN(n_0_0_182));
   OAI22_X1 i_0_0_360 (.A1(n_0_0_350), .A2(n_0_0_287), .B1(n_0_0_343), .B2(
      n_0_0_238), .ZN(n_0_0_183));
   INV_X1 i_0_0_361 (.A(n_0_0_185), .ZN(n_0_0_184));
   NAND2_X1 i_0_0_362 (.A1(n_0_0_187), .A2(n_0_0_186), .ZN(n_0_0_185));
   AOI22_X1 i_0_0_363 (.A1(op1[13]), .A2(n_0_0_305), .B1(op1[12]), .B2(n_0_0_303), 
      .ZN(n_0_0_186));
   AOI22_X1 i_0_0_364 (.A1(OP1_complement[13]), .A2(n_0_0_304), .B1(
      OP1_complement[12]), .B2(n_0_0_302), .ZN(n_0_0_187));
   OAI22_X1 i_0_0_365 (.A1(n[0]), .A2(n_0_0_201), .B1(n_0_0_356), .B2(n_0_0_188), 
      .ZN(n_0_134));
   AOI22_X1 i_0_0_366 (.A1(n[1]), .A2(n_0_0_189), .B1(n_0_0_357), .B2(n_0_0_215), 
      .ZN(n_0_0_188));
   AOI211_X1 i_0_0_367 (.A(n_0_0_194), .B(n_0_0_190), .C1(n_0_0_349), .C2(
      n_0_0_292), .ZN(n_0_0_189));
   OAI22_X1 i_0_0_368 (.A1(n_0_0_343), .A2(n_0_0_246), .B1(n_0_0_345), .B2(
      n_0_0_191), .ZN(n_0_0_190));
   NAND2_X1 i_0_0_369 (.A1(n_0_0_193), .A2(n_0_0_192), .ZN(n_0_0_191));
   AOI22_X1 i_0_0_370 (.A1(op1[14]), .A2(n_0_0_305), .B1(op1[13]), .B2(n_0_0_303), 
      .ZN(n_0_0_192));
   AOI22_X1 i_0_0_371 (.A1(OP1_complement[14]), .A2(n_0_0_304), .B1(
      OP1_complement[13]), .B2(n_0_0_302), .ZN(n_0_0_193));
   NOR2_X1 i_0_0_372 (.A1(n_0_0_340), .A2(n_0_89), .ZN(n_0_0_194));
   OAI22_X1 i_0_0_373 (.A1(n_0_0_356), .A2(n_0_0_195), .B1(n[0]), .B2(n_0_0_207), 
      .ZN(n_0_135));
   AOI22_X1 i_0_0_374 (.A1(n_0_0_357), .A2(n_0_0_222), .B1(n[1]), .B2(n_0_0_196), 
      .ZN(n_0_0_195));
   OAI21_X1 i_0_0_375 (.A(n_0_0_197), .B1(n_0_0_343), .B2(n_0_0_251), .ZN(
      n_0_0_196));
   AOI21_X1 i_0_0_376 (.A(n_0_0_244), .B1(n_0_0_344), .B2(n_0_0_198), .ZN(
      n_0_0_197));
   NAND2_X1 i_0_0_377 (.A1(n_0_0_200), .A2(n_0_0_199), .ZN(n_0_0_198));
   AOI22_X1 i_0_0_378 (.A1(op1[15]), .A2(n_0_0_305), .B1(op1[14]), .B2(n_0_0_303), 
      .ZN(n_0_0_199));
   AOI22_X1 i_0_0_379 (.A1(OP1_complement[15]), .A2(n_0_0_304), .B1(
      OP1_complement[14]), .B2(n_0_0_302), .ZN(n_0_0_200));
   OAI22_X1 i_0_0_380 (.A1(n_0_0_356), .A2(n_0_0_201), .B1(n[0]), .B2(n_0_0_214), 
      .ZN(n_0_136));
   AOI22_X1 i_0_0_381 (.A1(n_0_0_357), .A2(n_0_0_229), .B1(n[1]), .B2(n_0_0_202), 
      .ZN(n_0_0_201));
   OAI21_X1 i_0_0_382 (.A(n_0_0_203), .B1(n_0_0_343), .B2(n_0_0_257), .ZN(
      n_0_0_202));
   AOI21_X1 i_0_0_383 (.A(n_0_0_244), .B1(n_0_0_344), .B2(n_0_0_204), .ZN(
      n_0_0_203));
   NAND2_X1 i_0_0_384 (.A1(n_0_0_206), .A2(n_0_0_205), .ZN(n_0_0_204));
   AOI22_X1 i_0_0_385 (.A1(op1[16]), .A2(n_0_0_305), .B1(op1[15]), .B2(n_0_0_303), 
      .ZN(n_0_0_205));
   AOI22_X1 i_0_0_386 (.A1(OP1_complement[16]), .A2(n_0_0_304), .B1(
      OP1_complement[15]), .B2(n_0_0_302), .ZN(n_0_0_206));
   OAI22_X1 i_0_0_387 (.A1(n_0_0_356), .A2(n_0_0_207), .B1(n[0]), .B2(n_0_0_221), 
      .ZN(n_0_137));
   AOI22_X1 i_0_0_388 (.A1(n[1]), .A2(n_0_0_208), .B1(n_0_0_357), .B2(n_0_0_236), 
      .ZN(n_0_0_207));
   OAI21_X1 i_0_0_389 (.A(n_0_0_209), .B1(n_0_0_345), .B2(n_0_0_210), .ZN(
      n_0_0_208));
   AOI21_X1 i_0_0_390 (.A(n_0_0_244), .B1(n_0_0_342), .B2(n_0_0_263), .ZN(
      n_0_0_209));
   INV_X1 i_0_0_391 (.A(n_0_0_211), .ZN(n_0_0_210));
   NAND2_X1 i_0_0_392 (.A1(n_0_0_213), .A2(n_0_0_212), .ZN(n_0_0_211));
   AOI22_X1 i_0_0_393 (.A1(OP1_complement[17]), .A2(n_0_0_304), .B1(
      OP1_complement[16]), .B2(n_0_0_302), .ZN(n_0_0_212));
   AOI22_X1 i_0_0_394 (.A1(op1[17]), .A2(n_0_0_305), .B1(op1[16]), .B2(n_0_0_303), 
      .ZN(n_0_0_213));
   OAI22_X1 i_0_0_395 (.A1(n_0_0_356), .A2(n_0_0_214), .B1(n[0]), .B2(n_0_0_228), 
      .ZN(n_0_138));
   AOI22_X1 i_0_0_396 (.A1(n_0_0_357), .A2(n_0_0_242), .B1(n[1]), .B2(n_0_0_215), 
      .ZN(n_0_0_214));
   OAI21_X1 i_0_0_397 (.A(n_0_0_216), .B1(n_0_0_345), .B2(n_0_0_217), .ZN(
      n_0_0_215));
   AOI21_X1 i_0_0_398 (.A(n_0_0_244), .B1(n_0_0_342), .B2(n_0_0_269), .ZN(
      n_0_0_216));
   INV_X1 i_0_0_399 (.A(n_0_0_218), .ZN(n_0_0_217));
   NAND2_X1 i_0_0_400 (.A1(n_0_0_220), .A2(n_0_0_219), .ZN(n_0_0_218));
   AOI22_X1 i_0_0_401 (.A1(op1[18]), .A2(n_0_0_305), .B1(op1[17]), .B2(n_0_0_303), 
      .ZN(n_0_0_219));
   AOI22_X1 i_0_0_402 (.A1(OP1_complement[18]), .A2(n_0_0_304), .B1(
      OP1_complement[17]), .B2(n_0_0_302), .ZN(n_0_0_220));
   OAI22_X1 i_0_0_403 (.A1(n_0_0_356), .A2(n_0_0_221), .B1(n[0]), .B2(n_0_0_235), 
      .ZN(n_0_139));
   AOI22_X1 i_0_0_404 (.A1(n[1]), .A2(n_0_0_222), .B1(n_0_0_357), .B2(n_0_0_250), 
      .ZN(n_0_0_221));
   OAI21_X1 i_0_0_405 (.A(n_0_0_223), .B1(n_0_0_345), .B2(n_0_0_224), .ZN(
      n_0_0_222));
   AOI21_X1 i_0_0_406 (.A(n_0_0_244), .B1(n_0_0_342), .B2(n_0_0_275), .ZN(
      n_0_0_223));
   INV_X1 i_0_0_407 (.A(n_0_0_225), .ZN(n_0_0_224));
   NAND2_X1 i_0_0_408 (.A1(n_0_0_227), .A2(n_0_0_226), .ZN(n_0_0_225));
   AOI22_X1 i_0_0_409 (.A1(OP1_complement[19]), .A2(n_0_0_304), .B1(op1[18]), 
      .B2(n_0_0_303), .ZN(n_0_0_226));
   AOI22_X1 i_0_0_410 (.A1(op1[19]), .A2(n_0_0_305), .B1(OP1_complement[18]), 
      .B2(n_0_0_302), .ZN(n_0_0_227));
   OAI22_X1 i_0_0_411 (.A1(n_0_0_356), .A2(n_0_0_228), .B1(n[0]), .B2(n_0_0_241), 
      .ZN(n_0_140));
   AOI22_X1 i_0_0_412 (.A1(n[1]), .A2(n_0_0_229), .B1(n_0_0_357), .B2(n_0_0_256), 
      .ZN(n_0_0_228));
   OAI21_X1 i_0_0_413 (.A(n_0_0_230), .B1(n_0_0_345), .B2(n_0_0_231), .ZN(
      n_0_0_229));
   AOI21_X1 i_0_0_414 (.A(n_0_0_244), .B1(n_0_0_342), .B2(n_0_0_281), .ZN(
      n_0_0_230));
   INV_X1 i_0_0_415 (.A(n_0_0_232), .ZN(n_0_0_231));
   NAND2_X1 i_0_0_416 (.A1(n_0_0_234), .A2(n_0_0_233), .ZN(n_0_0_232));
   AOI22_X1 i_0_0_417 (.A1(op1[20]), .A2(n_0_0_305), .B1(op1[19]), .B2(n_0_0_303), 
      .ZN(n_0_0_233));
   AOI22_X1 i_0_0_418 (.A1(OP1_complement[20]), .A2(n_0_0_304), .B1(
      OP1_complement[19]), .B2(n_0_0_302), .ZN(n_0_0_234));
   OAI22_X1 i_0_0_419 (.A1(n_0_0_356), .A2(n_0_0_235), .B1(n[0]), .B2(n_0_0_249), 
      .ZN(n_0_141));
   AOI22_X1 i_0_0_420 (.A1(n[1]), .A2(n_0_0_236), .B1(n_0_0_357), .B2(n_0_0_261), 
      .ZN(n_0_0_235));
   OAI21_X1 i_0_0_421 (.A(n_0_0_237), .B1(n_0_0_343), .B2(n_0_0_286), .ZN(
      n_0_0_236));
   AOI21_X1 i_0_0_422 (.A(n_0_0_244), .B1(n_0_0_344), .B2(n_0_0_238), .ZN(
      n_0_0_237));
   NAND2_X1 i_0_0_423 (.A1(n_0_0_240), .A2(n_0_0_239), .ZN(n_0_0_238));
   AOI22_X1 i_0_0_424 (.A1(OP1_complement[21]), .A2(n_0_0_304), .B1(op1[20]), 
      .B2(n_0_0_303), .ZN(n_0_0_239));
   AOI22_X1 i_0_0_425 (.A1(op1[21]), .A2(n_0_0_305), .B1(OP1_complement[20]), 
      .B2(n_0_0_302), .ZN(n_0_0_240));
   OAI22_X1 i_0_0_426 (.A1(n_0_0_356), .A2(n_0_0_241), .B1(n[0]), .B2(n_0_0_255), 
      .ZN(n_0_142));
   AOI22_X1 i_0_0_427 (.A1(n[1]), .A2(n_0_0_242), .B1(n_0_0_357), .B2(n_0_0_267), 
      .ZN(n_0_0_241));
   OAI21_X1 i_0_0_428 (.A(n_0_0_243), .B1(n_0_0_345), .B2(n_0_0_245), .ZN(
      n_0_0_242));
   AOI21_X1 i_0_0_429 (.A(n_0_0_244), .B1(n_0_0_342), .B2(n_0_0_293), .ZN(
      n_0_0_243));
   NOR2_X1 i_0_0_430 (.A1(n[3]), .A2(n_0_0_299), .ZN(n_0_0_244));
   INV_X1 i_0_0_431 (.A(n_0_0_246), .ZN(n_0_0_245));
   NAND2_X1 i_0_0_432 (.A1(n_0_0_248), .A2(n_0_0_247), .ZN(n_0_0_246));
   AOI22_X1 i_0_0_433 (.A1(OP1_complement[22]), .A2(n_0_0_304), .B1(op1[21]), 
      .B2(n_0_0_303), .ZN(n_0_0_247));
   AOI22_X1 i_0_0_434 (.A1(op1[22]), .A2(n_0_0_305), .B1(OP1_complement[21]), 
      .B2(n_0_0_302), .ZN(n_0_0_248));
   OAI22_X1 i_0_0_435 (.A1(n_0_0_356), .A2(n_0_0_249), .B1(n[0]), .B2(n_0_0_260), 
      .ZN(n_0_143));
   AOI22_X1 i_0_0_436 (.A1(n_0_0_357), .A2(n_0_0_273), .B1(n[1]), .B2(n_0_0_250), 
      .ZN(n_0_0_249));
   AOI21_X1 i_0_0_437 (.A(n_0_0_296), .B1(n_0_0_344), .B2(n_0_0_251), .ZN(
      n_0_0_250));
   INV_X1 i_0_0_438 (.A(n_0_0_252), .ZN(n_0_0_251));
   NAND2_X1 i_0_0_439 (.A1(n_0_0_254), .A2(n_0_0_253), .ZN(n_0_0_252));
   AOI22_X1 i_0_0_440 (.A1(OP1_complement[23]), .A2(n_0_0_304), .B1(
      OP1_complement[22]), .B2(n_0_0_302), .ZN(n_0_0_253));
   AOI22_X1 i_0_0_441 (.A1(op1[23]), .A2(n_0_0_305), .B1(op1[22]), .B2(n_0_0_303), 
      .ZN(n_0_0_254));
   OAI22_X1 i_0_0_442 (.A1(n_0_0_356), .A2(n_0_0_255), .B1(n[0]), .B2(n_0_0_266), 
      .ZN(n_0_144));
   AOI22_X1 i_0_0_443 (.A1(n[1]), .A2(n_0_0_256), .B1(n_0_0_357), .B2(n_0_0_279), 
      .ZN(n_0_0_255));
   AOI21_X1 i_0_0_444 (.A(n_0_0_296), .B1(n_0_0_344), .B2(n_0_0_257), .ZN(
      n_0_0_256));
   AOI221_X1 i_0_0_445 (.A(n_0_0_258), .B1(op1[23]), .B2(n_0_0_303), .C1(
      OP1_complement[23]), .C2(n_0_0_302), .ZN(n_0_0_257));
   INV_X1 i_0_0_446 (.A(n_0_0_259), .ZN(n_0_0_258));
   AOI22_X1 i_0_0_447 (.A1(op1[24]), .A2(n_0_0_305), .B1(OP1_complement[24]), 
      .B2(n_0_0_304), .ZN(n_0_0_259));
   OAI22_X1 i_0_0_448 (.A1(n_0_0_356), .A2(n_0_0_260), .B1(n[0]), .B2(n_0_0_272), 
      .ZN(n_0_145));
   AOI22_X1 i_0_0_449 (.A1(n_0_0_357), .A2(n_0_0_285), .B1(n[1]), .B2(n_0_0_261), 
      .ZN(n_0_0_260));
   AOI21_X1 i_0_0_450 (.A(n_0_0_296), .B1(n_0_0_344), .B2(n_0_0_262), .ZN(
      n_0_0_261));
   INV_X1 i_0_0_451 (.A(n_0_0_263), .ZN(n_0_0_262));
   NAND2_X1 i_0_0_452 (.A1(n_0_0_265), .A2(n_0_0_264), .ZN(n_0_0_263));
   AOI22_X1 i_0_0_453 (.A1(OP1_complement[25]), .A2(n_0_0_304), .B1(op1[24]), 
      .B2(n_0_0_303), .ZN(n_0_0_264));
   AOI22_X1 i_0_0_454 (.A1(op1[25]), .A2(n_0_0_305), .B1(OP1_complement[24]), 
      .B2(n_0_0_302), .ZN(n_0_0_265));
   OAI22_X1 i_0_0_455 (.A1(n_0_0_356), .A2(n_0_0_266), .B1(n[0]), .B2(n_0_0_278), 
      .ZN(n_0_146));
   AOI22_X1 i_0_0_456 (.A1(n_0_0_357), .A2(n_0_0_291), .B1(n[1]), .B2(n_0_0_267), 
      .ZN(n_0_0_266));
   AOI21_X1 i_0_0_457 (.A(n_0_0_296), .B1(n_0_0_344), .B2(n_0_0_268), .ZN(
      n_0_0_267));
   INV_X1 i_0_0_458 (.A(n_0_0_269), .ZN(n_0_0_268));
   NAND2_X1 i_0_0_459 (.A1(n_0_0_271), .A2(n_0_0_270), .ZN(n_0_0_269));
   AOI22_X1 i_0_0_460 (.A1(OP1_complement[26]), .A2(n_0_0_304), .B1(
      OP1_complement[25]), .B2(n_0_0_302), .ZN(n_0_0_270));
   AOI22_X1 i_0_0_461 (.A1(op1[26]), .A2(n_0_0_305), .B1(op1[25]), .B2(n_0_0_303), 
      .ZN(n_0_0_271));
   OAI22_X1 i_0_0_462 (.A1(n_0_0_356), .A2(n_0_0_272), .B1(n[0]), .B2(n_0_0_284), 
      .ZN(n_0_147));
   AOI21_X1 i_0_0_463 (.A(n_0_0_297), .B1(n[1]), .B2(n_0_0_273), .ZN(n_0_0_272));
   AOI21_X1 i_0_0_464 (.A(n_0_0_296), .B1(n_0_0_344), .B2(n_0_0_274), .ZN(
      n_0_0_273));
   INV_X1 i_0_0_465 (.A(n_0_0_275), .ZN(n_0_0_274));
   NAND2_X1 i_0_0_466 (.A1(n_0_0_277), .A2(n_0_0_276), .ZN(n_0_0_275));
   AOI22_X1 i_0_0_467 (.A1(OP1_complement[27]), .A2(n_0_0_304), .B1(
      OP1_complement[26]), .B2(n_0_0_302), .ZN(n_0_0_276));
   AOI22_X1 i_0_0_468 (.A1(op1[27]), .A2(n_0_0_305), .B1(op1[26]), .B2(n_0_0_303), 
      .ZN(n_0_0_277));
   OAI22_X1 i_0_0_469 (.A1(n_0_0_356), .A2(n_0_0_278), .B1(n[0]), .B2(n_0_0_290), 
      .ZN(n_0_148));
   AOI21_X1 i_0_0_470 (.A(n_0_0_297), .B1(n[1]), .B2(n_0_0_279), .ZN(n_0_0_278));
   AOI21_X1 i_0_0_471 (.A(n_0_0_296), .B1(n_0_0_344), .B2(n_0_0_280), .ZN(
      n_0_0_279));
   INV_X1 i_0_0_472 (.A(n_0_0_281), .ZN(n_0_0_280));
   NAND2_X1 i_0_0_473 (.A1(n_0_0_283), .A2(n_0_0_282), .ZN(n_0_0_281));
   AOI22_X1 i_0_0_474 (.A1(OP1_complement[28]), .A2(n_0_0_304), .B1(op1[27]), 
      .B2(n_0_0_303), .ZN(n_0_0_282));
   AOI22_X1 i_0_0_475 (.A1(op1[28]), .A2(n_0_0_305), .B1(OP1_complement[27]), 
      .B2(n_0_0_302), .ZN(n_0_0_283));
   AOI21_X1 i_0_0_476 (.A(n_0_0_298), .B1(n[0]), .B2(n_0_0_284), .ZN(n_0_149));
   AOI21_X1 i_0_0_477 (.A(n_0_0_297), .B1(n[1]), .B2(n_0_0_285), .ZN(n_0_0_284));
   AOI21_X1 i_0_0_478 (.A(n_0_0_296), .B1(n_0_0_344), .B2(n_0_0_286), .ZN(
      n_0_0_285));
   INV_X1 i_0_0_479 (.A(n_0_0_287), .ZN(n_0_0_286));
   NAND2_X1 i_0_0_480 (.A1(n_0_0_289), .A2(n_0_0_288), .ZN(n_0_0_287));
   AOI22_X1 i_0_0_481 (.A1(op1[29]), .A2(n_0_0_305), .B1(OP1_complement[28]), 
      .B2(n_0_0_302), .ZN(n_0_0_288));
   AOI22_X1 i_0_0_482 (.A1(OP1_complement[29]), .A2(n_0_0_304), .B1(op1[28]), 
      .B2(n_0_0_303), .ZN(n_0_0_289));
   AOI21_X1 i_0_0_483 (.A(n_0_0_298), .B1(n[0]), .B2(n_0_0_290), .ZN(n_0_150));
   AOI21_X1 i_0_0_484 (.A(n_0_0_297), .B1(n[1]), .B2(n_0_0_291), .ZN(n_0_0_290));
   AOI21_X1 i_0_0_485 (.A(n_0_0_296), .B1(n_0_0_344), .B2(n_0_0_292), .ZN(
      n_0_0_291));
   INV_X1 i_0_0_486 (.A(n_0_0_293), .ZN(n_0_0_292));
   NAND2_X1 i_0_0_487 (.A1(n_0_0_295), .A2(n_0_0_294), .ZN(n_0_0_293));
   AOI22_X1 i_0_0_488 (.A1(OP1_complement[30]), .A2(n_0_0_304), .B1(
      OP1_complement[29]), .B2(n_0_0_302), .ZN(n_0_0_294));
   AOI22_X1 i_0_0_489 (.A1(op1[30]), .A2(n_0_0_305), .B1(op1[29]), .B2(n_0_0_303), 
      .ZN(n_0_0_295));
   NOR2_X1 i_0_0_490 (.A1(n_0_0_344), .A2(n_0_89), .ZN(n_0_0_296));
   NOR2_X1 i_0_0_491 (.A1(n[1]), .A2(n_0_0_299), .ZN(n_0_0_297));
   NOR2_X1 i_0_0_492 (.A1(n[0]), .A2(n_0_89), .ZN(n_0_0_298));
   INV_X1 i_0_0_493 (.A(n_0_89), .ZN(n_0_0_299));
   NAND2_X1 i_0_0_494 (.A1(n_0_0_301), .A2(n_0_0_300), .ZN(n_0_89));
   AOI22_X1 i_0_0_495 (.A1(OP1_complement[31]), .A2(n_0_0_304), .B1(op1[30]), 
      .B2(n_0_0_303), .ZN(n_0_0_300));
   AOI22_X1 i_0_0_496 (.A1(op1[31]), .A2(n_0_0_305), .B1(OP1_complement[30]), 
      .B2(n_0_0_302), .ZN(n_0_0_301));
   NOR3_X1 i_0_0_497 (.A1(q), .A2(n_0_0_327), .A3(n_0_0_306), .ZN(n_0_0_302));
   NOR3_X1 i_0_0_498 (.A1(n_0_0_355), .A2(n_0_0_326), .A3(n_0_0_307), .ZN(
      n_0_0_303));
   AND2_X1 i_0_0_499 (.A1(n_0_0_325), .A2(n_0_0_307), .ZN(n_0_0_304));
   AND2_X1 i_0_0_500 (.A1(n_0_0_325), .A2(n_0_0_306), .ZN(n_0_0_305));
   INV_X1 i_0_0_501 (.A(n_0_0_307), .ZN(n_0_0_306));
   NAND4_X1 i_0_0_502 (.A1(n_0_0_311), .A2(n_0_0_308), .A3(n_0_0_317), .A4(
      n_0_0_319), .ZN(n_0_0_307));
   AOI21_X1 i_0_0_503 (.A(n_0_0_309), .B1(op2[11]), .B2(n_0_0_348), .ZN(
      n_0_0_308));
   NOR3_X1 i_0_0_504 (.A1(n[0]), .A2(n_0_0_340), .A3(n_0_0_310), .ZN(n_0_0_309));
   AOI22_X1 i_0_0_505 (.A1(n_0_0_357), .A2(op2[1]), .B1(n[1]), .B2(op2[5]), 
      .ZN(n_0_0_310));
   AOI21_X1 i_0_0_506 (.A(n_0_0_312), .B1(op2[3]), .B2(n_0_0_338), .ZN(n_0_0_311));
   NOR3_X1 i_0_0_507 (.A1(n[0]), .A2(n_0_0_350), .A3(n_0_0_313), .ZN(n_0_0_312));
   AOI22_X1 i_0_0_508 (.A1(n_0_0_357), .A2(op2[9]), .B1(n[1]), .B2(op2[13]), 
      .ZN(n_0_0_313));
   INV_X1 i_0_0_509 (.A(n_0_0_315), .ZN(n_0_0_314));
   NAND2_X1 i_0_0_510 (.A1(n_0_0_358), .A2(n_0_0_316), .ZN(n_0_0_315));
   NOR2_X1 i_0_0_511 (.A1(n[3]), .A2(n[1]), .ZN(n_0_0_316));
   OR3_X1 i_0_0_512 (.A1(n_0_0_357), .A2(n_0_0_356), .A3(n_0_0_318), .ZN(
      n_0_0_317));
   AOI22_X1 i_0_0_513 (.A1(op2[15]), .A2(n_0_0_349), .B1(op2[7]), .B2(n_0_0_339), 
      .ZN(n_0_0_318));
   INV_X1 i_0_0_514 (.A(n_0_0_320), .ZN(n_0_0_319));
   OAI33_X1 i_0_0_515 (.A1(n_0_0_324), .A2(n_0_0_323), .A3(n_0_0_343), .B1(
      n_0_0_322), .B2(n_0_0_321), .B3(n_0_0_345), .ZN(n_0_0_320));
   AOI221_X1 i_0_0_516 (.A(n[1]), .B1(n_0_0_356), .B2(op2[25]), .C1(n[0]), 
      .C2(op2[27]), .ZN(n_0_0_321));
   AOI221_X1 i_0_0_517 (.A(n_0_0_357), .B1(n[0]), .B2(op2[31]), .C1(n_0_0_356), 
      .C2(op2[29]), .ZN(n_0_0_322));
   AOI221_X1 i_0_0_518 (.A(n_0_0_357), .B1(n[0]), .B2(op2[23]), .C1(n_0_0_356), 
      .C2(op2[21]), .ZN(n_0_0_323));
   AOI221_X1 i_0_0_519 (.A(n[1]), .B1(n_0_0_356), .B2(op2[17]), .C1(n[0]), 
      .C2(op2[19]), .ZN(n_0_0_324));
   AOI22_X1 i_0_0_520 (.A1(q), .A2(n_0_0_327), .B1(n_0_0_355), .B2(n_0_0_326), 
      .ZN(n_0_0_325));
   INV_X1 i_0_0_521 (.A(n_0_0_327), .ZN(n_0_0_326));
   NAND4_X1 i_0_0_522 (.A1(n_0_0_332), .A2(n_0_0_330), .A3(n_0_0_335), .A4(
      n_0_0_328), .ZN(n_0_0_327));
   INV_X1 i_0_0_523 (.A(n_0_0_329), .ZN(n_0_0_328));
   OAI33_X1 i_0_0_524 (.A1(n_0_0_346), .A2(n_0_0_345), .A3(n_0_0_357), .B1(n[1]), 
      .B2(n_0_0_356), .B3(n_0_0_341), .ZN(n_0_0_329));
   AOI221_X1 i_0_0_525 (.A(n_0_0_331), .B1(op2[10]), .B2(n_0_0_348), .C1(op2[2]), 
      .C2(n_0_0_338), .ZN(n_0_0_330));
   OAI33_X1 i_0_0_526 (.A1(n[0]), .A2(n_0_0_350), .A3(n_0_0_347), .B1(n[0]), 
      .B2(n_0_0_340), .B3(n_0_0_337), .ZN(n_0_0_331));
   OR3_X1 i_0_0_527 (.A1(n[0]), .A2(n_0_0_334), .A3(n_0_0_333), .ZN(n_0_0_332));
   AOI221_X1 i_0_0_528 (.A(n[1]), .B1(op2[24]), .B2(n_0_0_344), .C1(op2[16]), 
      .C2(n_0_0_342), .ZN(n_0_0_333));
   AOI21_X1 i_0_0_529 (.A(n_0_0_357), .B1(op2[20]), .B2(n_0_0_342), .ZN(
      n_0_0_334));
   OR3_X1 i_0_0_530 (.A1(n_0_0_357), .A2(n_0_0_356), .A3(n_0_0_336), .ZN(
      n_0_0_335));
   AOI222_X1 i_0_0_531 (.A1(op2[6]), .A2(n_0_0_339), .B1(op2[22]), .B2(n_0_0_342), 
      .C1(op2[14]), .C2(n_0_0_349), .ZN(n_0_0_336));
   AOI22_X1 i_0_0_532 (.A1(n_0_0_357), .A2(op2[0]), .B1(n[1]), .B2(op2[4]), 
      .ZN(n_0_0_337));
   NOR3_X1 i_0_0_533 (.A1(n[1]), .A2(n_0_0_356), .A3(n_0_0_340), .ZN(n_0_0_338));
   INV_X1 i_0_0_534 (.A(n_0_0_340), .ZN(n_0_0_339));
   NAND2_X1 i_0_0_535 (.A1(n_0_0_359), .A2(n_0_0_358), .ZN(n_0_0_340));
   AOI22_X1 i_0_0_536 (.A1(op2[26]), .A2(n_0_0_344), .B1(op2[18]), .B2(n_0_0_342), 
      .ZN(n_0_0_341));
   INV_X1 i_0_0_537 (.A(n_0_0_343), .ZN(n_0_0_342));
   NAND2_X1 i_0_0_538 (.A1(n[3]), .A2(n_0_0_358), .ZN(n_0_0_343));
   INV_X1 i_0_0_539 (.A(n_0_0_345), .ZN(n_0_0_344));
   NAND2_X1 i_0_0_540 (.A1(n[3]), .A2(n[2]), .ZN(n_0_0_345));
   AOI22_X1 i_0_0_541 (.A1(n_0_0_356), .A2(op2[28]), .B1(n[0]), .B2(op2[30]), 
      .ZN(n_0_0_346));
   AOI22_X1 i_0_0_542 (.A1(n_0_0_357), .A2(op2[8]), .B1(n[1]), .B2(op2[12]), 
      .ZN(n_0_0_347));
   NOR3_X1 i_0_0_543 (.A1(n[1]), .A2(n_0_0_356), .A3(n_0_0_350), .ZN(n_0_0_348));
   INV_X1 i_0_0_544 (.A(n_0_0_350), .ZN(n_0_0_349));
   NAND2_X1 i_0_0_545 (.A1(n_0_0_359), .A2(n[2]), .ZN(n_0_0_350));
   INV_X1 i_0_0_546 (.A(n_0_0_6), .ZN(n_0_0_351));
   INV_X1 i_0_0_547 (.A(n_0_0_5), .ZN(n_0_0_352));
   INV_X1 i_0_0_548 (.A(n_0_0_4), .ZN(n_0_0_353));
   INV_X1 i_0_0_549 (.A(rst), .ZN(n_0_0_354));
   INV_X1 i_0_0_550 (.A(q), .ZN(n_0_0_355));
   INV_X1 i_0_0_551 (.A(n[0]), .ZN(n_0_0_356));
   INV_X1 i_0_0_552 (.A(n[1]), .ZN(n_0_0_357));
   INV_X1 i_0_0_553 (.A(n[2]), .ZN(n_0_0_358));
   INV_X1 i_0_0_554 (.A(n[3]), .ZN(n_0_0_359));
   DFF_X1 \adder_reg[63]  (.D(n_0_278), .CK(n_0_88), .Q(adder[63]), .QN());
   DFF_X1 \adder_reg[62]  (.D(n_0_277), .CK(n_0_88), .Q(adder[62]), .QN());
   DFF_X1 \adder_reg[61]  (.D(n_0_276), .CK(n_0_88), .Q(adder[61]), .QN());
   DFF_X1 \adder_reg[60]  (.D(n_0_275), .CK(n_0_88), .Q(adder[60]), .QN());
   DFF_X1 \adder_reg[59]  (.D(n_0_274), .CK(n_0_88), .Q(adder[59]), .QN());
   DFF_X1 \adder_reg[58]  (.D(n_0_273), .CK(n_0_88), .Q(adder[58]), .QN());
   DFF_X1 \adder_reg[57]  (.D(n_0_272), .CK(n_0_88), .Q(adder[57]), .QN());
   DFF_X1 \adder_reg[56]  (.D(n_0_271), .CK(n_0_88), .Q(adder[56]), .QN());
   DFF_X1 \adder_reg[55]  (.D(n_0_270), .CK(n_0_88), .Q(adder[55]), .QN());
   DFF_X1 \adder_reg[54]  (.D(n_0_269), .CK(n_0_88), .Q(adder[54]), .QN());
   DFF_X1 \adder_reg[53]  (.D(n_0_268), .CK(n_0_88), .Q(adder[53]), .QN());
   DFF_X1 \adder_reg[52]  (.D(n_0_267), .CK(n_0_88), .Q(adder[52]), .QN());
   DFF_X1 \adder_reg[51]  (.D(n_0_266), .CK(n_0_88), .Q(adder[51]), .QN());
   DFF_X1 \adder_reg[50]  (.D(n_0_265), .CK(n_0_88), .Q(adder[50]), .QN());
   DFF_X1 \adder_reg[49]  (.D(n_0_264), .CK(n_0_88), .Q(adder[49]), .QN());
   DFF_X1 \adder_reg[48]  (.D(n_0_263), .CK(n_0_88), .Q(adder[48]), .QN());
   DFF_X1 \adder_reg[47]  (.D(n_0_262), .CK(n_0_88), .Q(adder[47]), .QN());
   DFF_X1 \adder_reg[46]  (.D(n_0_261), .CK(n_0_88), .Q(adder[46]), .QN());
   DFF_X1 \adder_reg[45]  (.D(n_0_260), .CK(n_0_88), .Q(adder[45]), .QN());
   DFF_X1 \adder_reg[44]  (.D(n_0_259), .CK(n_0_88), .Q(adder[44]), .QN());
   DFF_X1 \adder_reg[43]  (.D(n_0_258), .CK(n_0_88), .Q(adder[43]), .QN());
   DFF_X1 \adder_reg[42]  (.D(n_0_257), .CK(n_0_88), .Q(adder[42]), .QN());
   DFF_X1 \adder_reg[41]  (.D(n_0_256), .CK(n_0_88), .Q(adder[41]), .QN());
   DFF_X1 \adder_reg[40]  (.D(n_0_255), .CK(n_0_88), .Q(adder[40]), .QN());
   DFF_X1 \adder_reg[39]  (.D(n_0_254), .CK(n_0_88), .Q(adder[39]), .QN());
   DFF_X1 \adder_reg[38]  (.D(n_0_253), .CK(n_0_88), .Q(adder[38]), .QN());
   DFF_X1 \adder_reg[37]  (.D(n_0_252), .CK(n_0_88), .Q(adder[37]), .QN());
   DFF_X1 \adder_reg[36]  (.D(n_0_251), .CK(n_0_88), .Q(adder[36]), .QN());
   DFF_X1 \adder_reg[35]  (.D(n_0_250), .CK(n_0_88), .Q(adder[35]), .QN());
   DFF_X1 \adder_reg[34]  (.D(n_0_249), .CK(n_0_88), .Q(adder[34]), .QN());
   DFF_X1 \adder_reg[33]  (.D(n_0_248), .CK(n_0_88), .Q(adder[33]), .QN());
   DFF_X1 \adder_reg[32]  (.D(n_0_247), .CK(n_0_88), .Q(adder[32]), .QN());
   DFF_X1 \adder_reg[31]  (.D(n_0_246), .CK(n_0_88), .Q(adder[31]), .QN());
   DFF_X1 \adder_reg[30]  (.D(n_0_245), .CK(n_0_88), .Q(adder[30]), .QN());
   DFF_X1 \adder_reg[29]  (.D(n_0_244), .CK(n_0_88), .Q(adder[29]), .QN());
   DFF_X1 \adder_reg[28]  (.D(n_0_243), .CK(n_0_88), .Q(adder[28]), .QN());
   DFF_X1 \adder_reg[27]  (.D(n_0_242), .CK(n_0_88), .Q(adder[27]), .QN());
   DFF_X1 \adder_reg[26]  (.D(n_0_241), .CK(n_0_88), .Q(adder[26]), .QN());
   DFF_X1 \adder_reg[25]  (.D(n_0_240), .CK(n_0_88), .Q(adder[25]), .QN());
   DFF_X1 \adder_reg[24]  (.D(n_0_239), .CK(n_0_88), .Q(adder[24]), .QN());
   DFF_X1 \adder_reg[23]  (.D(n_0_238), .CK(n_0_88), .Q(adder[23]), .QN());
   DFF_X1 \adder_reg[22]  (.D(n_0_237), .CK(n_0_88), .Q(adder[22]), .QN());
   DFF_X1 \adder_reg[21]  (.D(n_0_236), .CK(n_0_88), .Q(adder[21]), .QN());
   DFF_X1 \adder_reg[20]  (.D(n_0_235), .CK(n_0_88), .Q(adder[20]), .QN());
   DFF_X1 \adder_reg[19]  (.D(n_0_234), .CK(n_0_88), .Q(adder[19]), .QN());
   DFF_X1 \adder_reg[18]  (.D(n_0_233), .CK(n_0_88), .Q(adder[18]), .QN());
   DFF_X1 \adder_reg[17]  (.D(n_0_232), .CK(n_0_88), .Q(adder[17]), .QN());
   DFF_X1 \adder_reg[16]  (.D(n_0_231), .CK(n_0_88), .Q(adder[16]), .QN());
   DFF_X1 \adder_reg[15]  (.D(n_0_230), .CK(n_0_88), .Q(adder[15]), .QN());
   DFF_X1 \adder_reg[14]  (.D(n_0_229), .CK(n_0_88), .Q(adder[14]), .QN());
   DFF_X1 \adder_reg[13]  (.D(n_0_228), .CK(n_0_88), .Q(adder[13]), .QN());
   DFF_X1 \adder_reg[12]  (.D(n_0_227), .CK(n_0_88), .Q(adder[12]), .QN());
   DFF_X1 \adder_reg[11]  (.D(n_0_226), .CK(n_0_88), .Q(adder[11]), .QN());
   DFF_X1 \adder_reg[10]  (.D(n_0_225), .CK(n_0_88), .Q(adder[10]), .QN());
   DFF_X1 \adder_reg[9]  (.D(n_0_224), .CK(n_0_88), .Q(adder[9]), .QN());
   DFF_X1 \adder_reg[8]  (.D(n_0_223), .CK(n_0_88), .Q(adder[8]), .QN());
   DFF_X1 \adder_reg[7]  (.D(n_0_222), .CK(n_0_88), .Q(adder[7]), .QN());
   DFF_X1 \adder_reg[6]  (.D(n_0_221), .CK(n_0_88), .Q(adder[6]), .QN());
   DFF_X1 \adder_reg[5]  (.D(n_0_220), .CK(n_0_88), .Q(adder[5]), .QN());
   DFF_X1 \adder_reg[4]  (.D(n_0_219), .CK(n_0_88), .Q(adder[4]), .QN());
   DFF_X1 \adder_reg[3]  (.D(n_0_218), .CK(n_0_88), .Q(adder[3]), .QN());
   DFF_X1 \adder_reg[2]  (.D(n_0_217), .CK(n_0_88), .Q(adder[2]), .QN());
   DFF_X1 \adder_reg[1]  (.D(n_0_216), .CK(n_0_88), .Q(adder[1]), .QN());
   DFF_X1 \adder_reg[0]  (.D(n_0_215), .CK(n_0_88), .Q(adder[0]), .QN());
   DFF_X1 \n_reg[5]  (.D(n_0_83), .CK(n_0_88), .Q(n[5]), .QN());
   DFF_X1 \n_reg[4]  (.D(n_0_82), .CK(n_0_88), .Q(n[4]), .QN());
   DFF_X1 \n_reg[3]  (.D(n_0_81), .CK(n_0_88), .Q(n[3]), .QN());
   DFF_X1 \n_reg[2]  (.D(n_0_80), .CK(n_0_88), .Q(n[2]), .QN());
   DFF_X1 \n_reg[1]  (.D(n_0_79), .CK(n_0_88), .Q(n[1]), .QN());
   DFF_X1 \n_reg[0]  (.D(n_0_78), .CK(n_0_88), .Q(n[0]), .QN());
   CLKGATETST_X1 clk_gate_OP1_complement_reg (.CK(clk), .E(rst), .SE(1'b0), 
      .GCK(n_0_87));
   DFF_X1 \OP1_complement_reg[31]  (.D(n_0_33), .CK(n_0_87), .Q(
      OP1_complement[31]), .QN());
   DFF_X1 \OP1_complement_reg[30]  (.D(n_0_32), .CK(n_0_87), .Q(
      OP1_complement[30]), .QN());
   DFF_X1 \OP1_complement_reg[29]  (.D(n_0_31), .CK(n_0_87), .Q(
      OP1_complement[29]), .QN());
   DFF_X1 \OP1_complement_reg[28]  (.D(n_0_30), .CK(n_0_87), .Q(
      OP1_complement[28]), .QN());
   DFF_X1 \OP1_complement_reg[27]  (.D(n_0_29), .CK(n_0_87), .Q(
      OP1_complement[27]), .QN());
   DFF_X1 \OP1_complement_reg[26]  (.D(n_0_28), .CK(n_0_87), .Q(
      OP1_complement[26]), .QN());
   DFF_X1 \OP1_complement_reg[25]  (.D(n_0_27), .CK(n_0_87), .Q(
      OP1_complement[25]), .QN());
   DFF_X1 \OP1_complement_reg[24]  (.D(n_0_26), .CK(n_0_87), .Q(
      OP1_complement[24]), .QN());
   DFF_X1 \OP1_complement_reg[23]  (.D(n_0_25), .CK(n_0_87), .Q(
      OP1_complement[23]), .QN());
   DFF_X1 \OP1_complement_reg[22]  (.D(n_0_24), .CK(n_0_87), .Q(
      OP1_complement[22]), .QN());
   DFF_X1 \OP1_complement_reg[21]  (.D(n_0_23), .CK(n_0_87), .Q(
      OP1_complement[21]), .QN());
   DFF_X1 \OP1_complement_reg[20]  (.D(n_0_22), .CK(n_0_87), .Q(
      OP1_complement[20]), .QN());
   DFF_X1 \OP1_complement_reg[19]  (.D(n_0_21), .CK(n_0_87), .Q(
      OP1_complement[19]), .QN());
   DFF_X1 \OP1_complement_reg[18]  (.D(n_0_20), .CK(n_0_87), .Q(
      OP1_complement[18]), .QN());
   DFF_X1 \OP1_complement_reg[17]  (.D(n_0_19), .CK(n_0_87), .Q(
      OP1_complement[17]), .QN());
   DFF_X1 \OP1_complement_reg[16]  (.D(n_0_18), .CK(n_0_87), .Q(
      OP1_complement[16]), .QN());
   DFF_X1 \OP1_complement_reg[15]  (.D(n_0_17), .CK(n_0_87), .Q(
      OP1_complement[15]), .QN());
   DFF_X1 \OP1_complement_reg[14]  (.D(n_0_16), .CK(n_0_87), .Q(
      OP1_complement[14]), .QN());
   DFF_X1 \OP1_complement_reg[13]  (.D(n_0_15), .CK(n_0_87), .Q(
      OP1_complement[13]), .QN());
   DFF_X1 \OP1_complement_reg[12]  (.D(n_0_14), .CK(n_0_87), .Q(
      OP1_complement[12]), .QN());
   DFF_X1 \OP1_complement_reg[11]  (.D(n_0_13), .CK(n_0_87), .Q(
      OP1_complement[11]), .QN());
   DFF_X1 \OP1_complement_reg[10]  (.D(n_0_12), .CK(n_0_87), .Q(
      OP1_complement[10]), .QN());
   DFF_X1 \OP1_complement_reg[9]  (.D(n_0_11), .CK(n_0_87), .Q(OP1_complement[9]), 
      .QN());
   DFF_X1 \OP1_complement_reg[8]  (.D(n_0_10), .CK(n_0_87), .Q(OP1_complement[8]), 
      .QN());
   DFF_X1 \OP1_complement_reg[7]  (.D(n_0_9), .CK(n_0_87), .Q(OP1_complement[7]), 
      .QN());
   DFF_X1 \OP1_complement_reg[6]  (.D(n_0_8), .CK(n_0_87), .Q(OP1_complement[6]), 
      .QN());
   DFF_X1 \OP1_complement_reg[5]  (.D(n_0_7), .CK(n_0_87), .Q(OP1_complement[5]), 
      .QN());
   DFF_X1 \OP1_complement_reg[4]  (.D(n_0_6), .CK(n_0_87), .Q(OP1_complement[4]), 
      .QN());
   DFF_X1 \OP1_complement_reg[3]  (.D(n_0_5), .CK(n_0_87), .Q(OP1_complement[3]), 
      .QN());
   DFF_X1 \OP1_complement_reg[2]  (.D(n_0_4), .CK(n_0_87), .Q(OP1_complement[2]), 
      .QN());
   DFF_X1 \OP1_complement_reg[1]  (.D(n_0_3), .CK(n_0_87), .Q(OP1_complement[1]), 
      .QN());
   DFF_X1 \OP1_complement_reg[0]  (.D(op1[0]), .CK(n_0_87), .Q(OP1_complement[0]), 
      .QN());
   DFF_X1 q_reg (.D(n_0_85), .CK(n_0_88), .Q(q), .QN());
   CLKGATETST_X1 clk_gate_adder_reg (.CK(clk), .E(n_0_84), .SE(1'b0), .GCK(
      n_0_88));
endmodule
