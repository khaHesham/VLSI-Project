
// 	Wed Jan  4 13:53:51 2023
//	vlsi
//	localhost.localdomain

module datapath__0_1 (M, A, p_0);

output [31:0] p_0;
input [31:0] A;
input [31:0] M;
wire n_0;
wire n_154;
wire n_1;
wire n_153;
wire n_152;
wire n_2;
wire n_157;
wire n_151;
wire n_3;
wire n_158;
wire n_164;
wire n_161;
wire n_149;
wire n_10;
wire n_9;
wire n_6;
wire n_7;
wire n_4;
wire n_146;
wire n_137;
wire n_11;
wire n_5;
wire n_147;
wire n_141;
wire n_8;
wire n_144;
wire n_142;
wire n_148;
wire n_139;
wire n_135;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_12;
wire n_132;
wire n_123;
wire n_19;
wire n_13;
wire n_133;
wire n_127;
wire n_16;
wire n_130;
wire n_128;
wire n_134;
wire n_125;
wire n_121;
wire n_26;
wire n_25;
wire n_22;
wire n_23;
wire n_20;
wire n_118;
wire n_109;
wire n_27;
wire n_21;
wire n_119;
wire n_113;
wire n_24;
wire n_116;
wire n_114;
wire n_120;
wire n_111;
wire n_107;
wire n_34;
wire n_33;
wire n_30;
wire n_31;
wire n_28;
wire n_104;
wire n_95;
wire n_35;
wire n_29;
wire n_105;
wire n_99;
wire n_32;
wire n_102;
wire n_100;
wire n_106;
wire n_97;
wire n_93;
wire n_42;
wire n_41;
wire n_38;
wire n_39;
wire n_36;
wire n_82;
wire n_72;
wire n_43;
wire n_37;
wire n_81;
wire n_84;
wire n_74;
wire n_40;
wire n_83;
wire n_79;
wire n_76;
wire n_86;
wire n_51;
wire n_50;
wire n_49;
wire n_47;
wire n_45;
wire n_44;
wire n_91;
wire n_48;
wire n_66;
wire n_53;
wire n_46;
wire n_90;
wire n_88;
wire n_69;
wire n_52;
wire n_71;
wire n_78;
wire n_165;
wire n_162;
wire n_64;
wire n_63;
wire n_62;
wire n_58;
wire n_55;
wire n_54;
wire n_160;
wire n_166;
wire n_163;
wire n_61;
wire n_60;
wire n_57;
wire n_56;
wire n_59;
wire n_159;
wire n_67;
wire n_65;
wire n_70;
wire n_77;
wire n_92;
wire n_89;
wire n_68;
wire n_87;
wire n_73;
wire n_85;
wire n_80;
wire n_75;
wire n_94;
wire n_98;
wire n_101;
wire n_96;
wire n_103;
wire n_108;
wire n_112;
wire n_115;
wire n_110;
wire n_117;
wire n_122;
wire n_126;
wire n_129;
wire n_124;
wire n_131;
wire n_136;
wire n_140;
wire n_143;
wire n_138;
wire n_145;
wire n_150;
wire n_156;
wire n_155;


INV_X1 i_198 (.ZN (n_166), .A (M[30]));
INV_X1 i_197 (.ZN (n_165), .A (M[27]));
INV_X1 i_196 (.ZN (n_164), .A (M[3]));
INV_X1 i_195 (.ZN (n_163), .A (A[31]));
INV_X1 i_194 (.ZN (n_162), .A (A[27]));
INV_X1 i_193 (.ZN (n_161), .A (A[3]));
NAND2_X1 i_192 (.ZN (n_160), .A1 (n_166), .A2 (n_163));
NOR2_X1 i_191 (.ZN (n_159), .A1 (M[28]), .A2 (A[28]));
NAND2_X1 i_190 (.ZN (n_158), .A1 (n_164), .A2 (n_161));
NAND2_X1 i_189 (.ZN (n_157), .A1 (M[2]), .A2 (A[2]));
INV_X1 i_188 (.ZN (n_156), .A (n_157));
NOR2_X1 i_187 (.ZN (n_155), .A1 (M[1]), .A2 (A[1]));
NAND2_X1 i_186 (.ZN (n_154), .A1 (M[0]), .A2 (A[0]));
NAND2_X1 i_185 (.ZN (n_153), .A1 (M[1]), .A2 (A[1]));
AOI21_X1 i_184 (.ZN (n_152), .A (n_155), .B1 (n_154), .B2 (n_153));
OAI22_X1 i_183 (.ZN (n_151), .A1 (M[2]), .A2 (A[2]), .B1 (n_156), .B2 (n_152));
OAI21_X1 i_182 (.ZN (n_150), .A (n_151), .B1 (n_164), .B2 (n_161));
NAND2_X1 i_181 (.ZN (n_149), .A1 (n_158), .A2 (n_150));
NOR2_X1 i_180 (.ZN (n_148), .A1 (M[7]), .A2 (A[7]));
NOR2_X1 i_179 (.ZN (n_147), .A1 (M[5]), .A2 (A[5]));
NOR2_X1 i_178 (.ZN (n_146), .A1 (M[6]), .A2 (A[6]));
OR3_X1 i_177 (.ZN (n_145), .A1 (n_148), .A2 (n_146), .A3 (n_147));
NOR2_X1 i_176 (.ZN (n_144), .A1 (M[4]), .A2 (A[4]));
NOR3_X1 i_175 (.ZN (n_143), .A1 (n_145), .A2 (n_144), .A3 (n_149));
NAND2_X1 i_174 (.ZN (n_142), .A1 (M[4]), .A2 (A[4]));
NAND2_X1 i_173 (.ZN (n_141), .A1 (M[5]), .A2 (A[5]));
AOI21_X1 i_172 (.ZN (n_140), .A (n_145), .B1 (n_142), .B2 (n_141));
AND2_X1 i_171 (.ZN (n_139), .A1 (M[7]), .A2 (A[7]));
NAND2_X1 i_170 (.ZN (n_138), .A1 (M[6]), .A2 (A[6]));
INV_X1 i_169 (.ZN (n_137), .A (n_138));
NOR2_X1 i_168 (.ZN (n_136), .A1 (n_148), .A2 (n_138));
NOR4_X1 i_167 (.ZN (n_135), .A1 (n_139), .A2 (n_136), .A3 (n_140), .A4 (n_143));
NOR2_X1 i_166 (.ZN (n_134), .A1 (M[11]), .A2 (A[11]));
NOR2_X1 i_165 (.ZN (n_133), .A1 (M[9]), .A2 (A[9]));
NOR2_X1 i_164 (.ZN (n_132), .A1 (M[10]), .A2 (A[10]));
OR3_X1 i_163 (.ZN (n_131), .A1 (n_134), .A2 (n_132), .A3 (n_133));
NOR2_X1 i_162 (.ZN (n_130), .A1 (M[8]), .A2 (A[8]));
NOR3_X1 i_161 (.ZN (n_129), .A1 (n_131), .A2 (n_130), .A3 (n_135));
NAND2_X1 i_160 (.ZN (n_128), .A1 (M[8]), .A2 (A[8]));
NAND2_X1 i_159 (.ZN (n_127), .A1 (M[9]), .A2 (A[9]));
AOI21_X1 i_158 (.ZN (n_126), .A (n_131), .B1 (n_128), .B2 (n_127));
AND2_X1 i_157 (.ZN (n_125), .A1 (M[11]), .A2 (A[11]));
NAND2_X1 i_156 (.ZN (n_124), .A1 (M[10]), .A2 (A[10]));
INV_X1 i_155 (.ZN (n_123), .A (n_124));
NOR2_X1 i_154 (.ZN (n_122), .A1 (n_134), .A2 (n_124));
NOR4_X1 i_153 (.ZN (n_121), .A1 (n_125), .A2 (n_122), .A3 (n_126), .A4 (n_129));
NOR2_X1 i_152 (.ZN (n_120), .A1 (M[15]), .A2 (A[15]));
NOR2_X1 i_151 (.ZN (n_119), .A1 (M[13]), .A2 (A[13]));
NOR2_X1 i_150 (.ZN (n_118), .A1 (M[14]), .A2 (A[14]));
OR3_X1 i_149 (.ZN (n_117), .A1 (n_120), .A2 (n_118), .A3 (n_119));
NOR2_X1 i_148 (.ZN (n_116), .A1 (M[12]), .A2 (A[12]));
NOR3_X1 i_147 (.ZN (n_115), .A1 (n_117), .A2 (n_116), .A3 (n_121));
NAND2_X1 i_146 (.ZN (n_114), .A1 (M[12]), .A2 (A[12]));
NAND2_X1 i_145 (.ZN (n_113), .A1 (M[13]), .A2 (A[13]));
AOI21_X1 i_144 (.ZN (n_112), .A (n_117), .B1 (n_114), .B2 (n_113));
AND2_X1 i_143 (.ZN (n_111), .A1 (M[15]), .A2 (A[15]));
NAND2_X1 i_142 (.ZN (n_110), .A1 (M[14]), .A2 (A[14]));
INV_X1 i_141 (.ZN (n_109), .A (n_110));
NOR2_X1 i_140 (.ZN (n_108), .A1 (n_120), .A2 (n_110));
NOR4_X1 i_139 (.ZN (n_107), .A1 (n_111), .A2 (n_108), .A3 (n_112), .A4 (n_115));
NOR2_X1 i_138 (.ZN (n_106), .A1 (M[19]), .A2 (A[19]));
NOR2_X1 i_137 (.ZN (n_105), .A1 (M[17]), .A2 (A[17]));
NOR2_X1 i_136 (.ZN (n_104), .A1 (M[18]), .A2 (A[18]));
OR3_X1 i_135 (.ZN (n_103), .A1 (n_106), .A2 (n_104), .A3 (n_105));
NOR2_X1 i_134 (.ZN (n_102), .A1 (M[16]), .A2 (A[16]));
NOR3_X1 i_133 (.ZN (n_101), .A1 (n_103), .A2 (n_102), .A3 (n_107));
NAND2_X1 i_132 (.ZN (n_100), .A1 (M[16]), .A2 (A[16]));
NAND2_X1 i_131 (.ZN (n_99), .A1 (M[17]), .A2 (A[17]));
AOI21_X1 i_130 (.ZN (n_98), .A (n_103), .B1 (n_100), .B2 (n_99));
AND2_X1 i_129 (.ZN (n_97), .A1 (M[19]), .A2 (A[19]));
NAND2_X1 i_128 (.ZN (n_96), .A1 (M[18]), .A2 (A[18]));
INV_X1 i_127 (.ZN (n_95), .A (n_96));
NOR2_X1 i_126 (.ZN (n_94), .A1 (n_106), .A2 (n_96));
NOR4_X1 i_125 (.ZN (n_93), .A1 (n_97), .A2 (n_94), .A3 (n_98), .A4 (n_101));
NOR2_X1 i_124 (.ZN (n_92), .A1 (M[27]), .A2 (A[27]));
NOR2_X1 i_123 (.ZN (n_91), .A1 (M[25]), .A2 (A[25]));
OAI22_X1 i_122 (.ZN (n_90), .A1 (M[25]), .A2 (A[25]), .B1 (M[26]), .B2 (A[26]));
OR2_X1 i_121 (.ZN (n_89), .A1 (n_92), .A2 (n_90));
NOR2_X1 i_120 (.ZN (n_88), .A1 (M[24]), .A2 (A[24]));
OR2_X1 i_119 (.ZN (n_87), .A1 (n_89), .A2 (n_88));
NOR2_X1 i_118 (.ZN (n_86), .A1 (M[23]), .A2 (A[23]));
INV_X1 i_117 (.ZN (n_85), .A (n_86));
NOR2_X1 i_116 (.ZN (n_84), .A1 (M[21]), .A2 (A[21]));
INV_X1 i_115 (.ZN (n_83), .A (n_84));
NOR2_X1 i_114 (.ZN (n_82), .A1 (M[22]), .A2 (A[22]));
INV_X1 i_113 (.ZN (n_81), .A (n_82));
NAND3_X1 i_112 (.ZN (n_80), .A1 (n_85), .A2 (n_81), .A3 (n_83));
NOR2_X1 i_111 (.ZN (n_79), .A1 (M[20]), .A2 (A[20]));
OR2_X1 i_110 (.ZN (n_78), .A1 (n_80), .A2 (n_79));
NOR3_X1 i_109 (.ZN (n_77), .A1 (n_87), .A2 (n_78), .A3 (n_93));
NAND2_X1 i_108 (.ZN (n_76), .A1 (M[20]), .A2 (A[20]));
NAND2_X1 i_107 (.ZN (n_75), .A1 (M[21]), .A2 (A[21]));
INV_X1 i_106 (.ZN (n_74), .A (n_75));
AOI21_X1 i_105 (.ZN (n_73), .A (n_80), .B1 (n_76), .B2 (n_75));
AND2_X1 i_104 (.ZN (n_72), .A1 (M[22]), .A2 (A[22]));
AOI221_X1 i_103 (.ZN (n_71), .A (n_73), .B1 (M[23]), .B2 (A[23]), .C1 (n_85), .C2 (n_72));
NOR2_X1 i_102 (.ZN (n_70), .A1 (n_87), .A2 (n_71));
NAND2_X1 i_101 (.ZN (n_69), .A1 (M[24]), .A2 (A[24]));
NAND2_X1 i_100 (.ZN (n_68), .A1 (M[25]), .A2 (A[25]));
AOI21_X1 i_99 (.ZN (n_67), .A (n_89), .B1 (n_69), .B2 (n_68));
NAND2_X1 i_98 (.ZN (n_66), .A1 (M[26]), .A2 (A[26]));
OAI22_X1 i_97 (.ZN (n_65), .A1 (n_165), .A2 (n_162), .B1 (n_92), .B2 (n_66));
NOR4_X1 i_96 (.ZN (n_64), .A1 (n_67), .A2 (n_65), .A3 (n_70), .A4 (n_77));
AOI21_X1 i_95 (.ZN (n_63), .A (n_159), .B1 (M[28]), .B2 (A[28]));
AOI21_X1 i_94 (.ZN (n_62), .A (n_159), .B1 (n_64), .B2 (n_63));
AOI21_X1 i_93 (.ZN (n_61), .A (n_62), .B1 (M[29]), .B2 (A[29]));
NOR2_X1 i_92 (.ZN (n_60), .A1 (M[29]), .A2 (A[29]));
OAI22_X1 i_91 (.ZN (n_59), .A1 (n_166), .A2 (n_163), .B1 (M[29]), .B2 (A[29]));
AOI21_X1 i_90 (.ZN (n_58), .A (n_60), .B1 (M[29]), .B2 (A[29]));
OAI21_X1 i_89 (.ZN (n_57), .A (n_160), .B1 (n_61), .B2 (n_59));
XNOR2_X1 i_88 (.ZN (n_56), .A (M[31]), .B (M[30]));
XOR2_X1 i_87 (.Z (p_0[31]), .A (n_57), .B (n_56));
NOR2_X1 i_86 (.ZN (n_55), .A1 (n_61), .A2 (n_60));
OAI21_X1 i_85 (.ZN (n_54), .A (n_160), .B1 (n_166), .B2 (n_163));
XNOR2_X1 i_84 (.ZN (p_0[30]), .A (n_55), .B (n_54));
XOR2_X1 i_83 (.Z (p_0[29]), .A (n_62), .B (n_58));
XNOR2_X1 i_82 (.ZN (p_0[28]), .A (n_64), .B (n_63));
OAI22_X1 i_81 (.ZN (n_53), .A1 (M[27]), .A2 (A[27]), .B1 (n_165), .B2 (n_162));
OAI21_X1 i_80 (.ZN (n_52), .A (n_71), .B1 (n_93), .B2 (n_78));
INV_X1 i_79 (.ZN (n_51), .A (n_52));
OAI21_X1 i_78 (.ZN (n_50), .A (n_69), .B1 (M[24]), .B2 (A[24]));
AOI21_X1 i_77 (.ZN (n_49), .A (n_88), .B1 (n_69), .B2 (n_51));
AOI21_X1 i_76 (.ZN (n_48), .A (n_49), .B1 (M[25]), .B2 (A[25]));
AOI21_X1 i_75 (.ZN (n_47), .A (n_91), .B1 (M[25]), .B2 (A[25]));
OAI21_X1 i_74 (.ZN (n_46), .A (n_66), .B1 (n_90), .B2 (n_48));
XNOR2_X1 i_73 (.ZN (p_0[27]), .A (n_53), .B (n_46));
OAI21_X1 i_72 (.ZN (n_45), .A (n_66), .B1 (M[26]), .B2 (A[26]));
NOR2_X1 i_71 (.ZN (n_44), .A1 (n_91), .A2 (n_48));
XNOR2_X1 i_70 (.ZN (p_0[26]), .A (n_45), .B (n_44));
XOR2_X1 i_69 (.Z (p_0[25]), .A (n_49), .B (n_47));
XOR2_X1 i_68 (.Z (p_0[24]), .A (n_51), .B (n_50));
AOI21_X1 i_67 (.ZN (n_43), .A (n_86), .B1 (M[23]), .B2 (A[23]));
OAI21_X1 i_66 (.ZN (n_42), .A (n_76), .B1 (M[20]), .B2 (A[20]));
AOI21_X1 i_65 (.ZN (n_41), .A (n_79), .B1 (n_93), .B2 (n_76));
OAI21_X1 i_64 (.ZN (n_40), .A (n_83), .B1 (n_74), .B2 (n_41));
INV_X1 i_63 (.ZN (n_39), .A (n_40));
NOR2_X1 i_62 (.ZN (n_38), .A1 (n_84), .A2 (n_74));
OAI21_X1 i_61 (.ZN (n_37), .A (n_81), .B1 (n_72), .B2 (n_39));
XNOR2_X1 i_60 (.ZN (p_0[23]), .A (n_43), .B (n_37));
NOR2_X1 i_59 (.ZN (n_36), .A1 (n_82), .A2 (n_72));
XOR2_X1 i_58 (.Z (p_0[22]), .A (n_39), .B (n_36));
XOR2_X1 i_57 (.Z (p_0[21]), .A (n_41), .B (n_38));
XOR2_X1 i_56 (.Z (p_0[20]), .A (n_93), .B (n_42));
NOR2_X1 i_55 (.ZN (n_35), .A1 (n_106), .A2 (n_97));
OAI21_X1 i_54 (.ZN (n_34), .A (n_100), .B1 (M[16]), .B2 (A[16]));
AOI21_X1 i_53 (.ZN (n_33), .A (n_102), .B1 (n_107), .B2 (n_100));
INV_X1 i_52 (.ZN (n_32), .A (n_33));
AOI21_X1 i_51 (.ZN (n_31), .A (n_105), .B1 (n_99), .B2 (n_32));
AOI21_X1 i_50 (.ZN (n_30), .A (n_105), .B1 (M[17]), .B2 (A[17]));
OAI22_X1 i_49 (.ZN (n_29), .A1 (M[18]), .A2 (A[18]), .B1 (n_95), .B2 (n_31));
XNOR2_X1 i_48 (.ZN (p_0[19]), .A (n_35), .B (n_29));
NOR2_X1 i_47 (.ZN (n_28), .A1 (n_104), .A2 (n_95));
XOR2_X1 i_46 (.Z (p_0[18]), .A (n_31), .B (n_28));
XOR2_X1 i_45 (.Z (p_0[17]), .A (n_33), .B (n_30));
XOR2_X1 i_44 (.Z (p_0[16]), .A (n_107), .B (n_34));
NOR2_X1 i_43 (.ZN (n_27), .A1 (n_120), .A2 (n_111));
OAI21_X1 i_42 (.ZN (n_26), .A (n_114), .B1 (M[12]), .B2 (A[12]));
AOI21_X1 i_41 (.ZN (n_25), .A (n_116), .B1 (n_121), .B2 (n_114));
INV_X1 i_40 (.ZN (n_24), .A (n_25));
AOI21_X1 i_39 (.ZN (n_23), .A (n_119), .B1 (n_113), .B2 (n_24));
AOI21_X1 i_38 (.ZN (n_22), .A (n_119), .B1 (M[13]), .B2 (A[13]));
OAI22_X1 i_37 (.ZN (n_21), .A1 (M[14]), .A2 (A[14]), .B1 (n_109), .B2 (n_23));
XNOR2_X1 i_36 (.ZN (p_0[15]), .A (n_27), .B (n_21));
NOR2_X1 i_35 (.ZN (n_20), .A1 (n_118), .A2 (n_109));
XOR2_X1 i_34 (.Z (p_0[14]), .A (n_23), .B (n_20));
XOR2_X1 i_33 (.Z (p_0[13]), .A (n_25), .B (n_22));
XOR2_X1 i_32 (.Z (p_0[12]), .A (n_121), .B (n_26));
NOR2_X1 i_31 (.ZN (n_19), .A1 (n_134), .A2 (n_125));
AOI21_X1 i_30 (.ZN (n_18), .A (n_130), .B1 (M[8]), .B2 (A[8]));
AOI21_X1 i_29 (.ZN (n_17), .A (n_130), .B1 (n_135), .B2 (n_128));
INV_X1 i_28 (.ZN (n_16), .A (n_17));
AOI21_X1 i_27 (.ZN (n_15), .A (n_133), .B1 (n_127), .B2 (n_16));
AOI21_X1 i_26 (.ZN (n_14), .A (n_133), .B1 (M[9]), .B2 (A[9]));
OAI22_X1 i_25 (.ZN (n_13), .A1 (M[10]), .A2 (A[10]), .B1 (n_123), .B2 (n_15));
XNOR2_X1 i_24 (.ZN (p_0[11]), .A (n_19), .B (n_13));
NOR2_X1 i_23 (.ZN (n_12), .A1 (n_132), .A2 (n_123));
XOR2_X1 i_22 (.Z (p_0[10]), .A (n_15), .B (n_12));
XOR2_X1 i_21 (.Z (p_0[9]), .A (n_17), .B (n_14));
XNOR2_X1 i_20 (.ZN (p_0[8]), .A (n_135), .B (n_18));
NOR2_X1 i_19 (.ZN (n_11), .A1 (n_148), .A2 (n_139));
OAI21_X1 i_18 (.ZN (n_10), .A (n_142), .B1 (M[4]), .B2 (A[4]));
AOI21_X1 i_17 (.ZN (n_9), .A (n_144), .B1 (n_149), .B2 (n_142));
INV_X1 i_16 (.ZN (n_8), .A (n_9));
AOI21_X1 i_15 (.ZN (n_7), .A (n_147), .B1 (n_141), .B2 (n_8));
AOI21_X1 i_14 (.ZN (n_6), .A (n_147), .B1 (M[5]), .B2 (A[5]));
OAI22_X1 i_13 (.ZN (n_5), .A1 (M[6]), .A2 (A[6]), .B1 (n_137), .B2 (n_7));
XNOR2_X1 i_12 (.ZN (p_0[7]), .A (n_11), .B (n_5));
NOR2_X1 i_11 (.ZN (n_4), .A1 (n_146), .A2 (n_137));
XOR2_X1 i_10 (.Z (p_0[6]), .A (n_7), .B (n_4));
XOR2_X1 i_9 (.Z (p_0[5]), .A (n_9), .B (n_6));
XOR2_X1 i_8 (.Z (p_0[4]), .A (n_149), .B (n_10));
OAI21_X1 i_7 (.ZN (n_3), .A (n_158), .B1 (n_164), .B2 (n_161));
XOR2_X1 i_6 (.Z (p_0[3]), .A (n_151), .B (n_3));
OAI21_X1 i_5 (.ZN (n_2), .A (n_157), .B1 (M[2]), .B2 (A[2]));
XNOR2_X1 i_4 (.ZN (p_0[2]), .A (n_152), .B (n_2));
OAI21_X1 i_3 (.ZN (n_1), .A (n_153), .B1 (M[1]), .B2 (A[1]));
XOR2_X1 i_2 (.Z (p_0[1]), .A (n_154), .B (n_1));
OAI21_X1 i_1 (.ZN (n_0), .A (n_154), .B1 (M[0]), .B2 (A[0]));
INV_X1 i_0 (.ZN (p_0[0]), .A (n_0));

endmodule //datapath__0_1

module datapath (A, p_0, M);

output [31:0] p_0;
input [31:0] A;
input [31:0] M;
wire n_0;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire n_12;
wire n_13;
wire n_14;
wire n_15;
wire n_16;
wire n_17;
wire n_18;
wire n_19;
wire n_20;
wire n_21;
wire n_22;
wire n_23;
wire n_24;
wire n_25;
wire n_26;
wire n_27;
wire n_28;
wire n_29;
wire n_30;
wire n_31;
wire n_32;
wire n_33;
wire n_34;
wire n_35;
wire n_36;
wire n_37;
wire n_38;
wire n_39;
wire n_40;
wire n_41;
wire n_42;
wire n_43;
wire n_44;
wire n_45;
wire n_46;
wire n_47;
wire n_48;
wire n_49;
wire n_50;
wire n_51;
wire n_52;
wire n_53;
wire n_54;
wire n_55;
wire n_56;
wire n_57;
wire n_58;
wire n_59;
wire n_60;
wire n_61;
wire n_62;
wire n_63;
wire n_64;
wire n_65;
wire n_66;
wire n_67;
wire n_68;
wire n_69;
wire n_70;
wire n_71;
wire n_72;
wire n_73;
wire n_74;
wire n_75;
wire n_76;
wire n_77;
wire n_78;
wire n_79;
wire n_80;
wire n_81;
wire n_82;
wire n_83;
wire n_84;
wire n_85;
wire n_86;
wire n_87;
wire n_88;
wire n_89;
wire n_90;
wire n_91;
wire n_92;
wire n_93;
wire n_94;


XNOR2_X1 i_126 (.ZN (p_0[31]), .A (n_94), .B (M[31]));
OAI33_X1 i_125 (.ZN (n_94), .A1 (n_93), .A2 (A[31]), .A3 (M[30]), .B1 (n_89), .B2 (n_90), .B3 (n_91));
INV_X1 i_124 (.ZN (n_93), .A (n_89));
XNOR2_X1 i_123 (.ZN (p_0[30]), .A (n_89), .B (n_92));
AOI22_X1 i_122 (.ZN (n_92), .A1 (n_90), .A2 (n_91), .B1 (A[31]), .B2 (M[30]));
INV_X1 i_121 (.ZN (n_91), .A (M[30]));
INV_X1 i_120 (.ZN (n_90), .A (A[31]));
AOI22_X1 i_119 (.ZN (n_89), .A1 (n_86), .A2 (n_87), .B1 (n_88), .B2 (M[29]));
INV_X1 i_118 (.ZN (n_88), .A (A[29]));
XNOR2_X1 i_117 (.ZN (p_0[29]), .A (n_86), .B (n_87));
XNOR2_X1 i_116 (.ZN (n_87), .A (A[29]), .B (M[29]));
OAI22_X1 i_115 (.ZN (n_86), .A1 (n_83), .A2 (n_84), .B1 (n_85), .B2 (A[28]));
INV_X1 i_114 (.ZN (n_85), .A (M[28]));
XNOR2_X1 i_113 (.ZN (p_0[28]), .A (n_83), .B (n_84));
XOR2_X1 i_112 (.Z (n_84), .A (A[28]), .B (M[28]));
AOI22_X1 i_111 (.ZN (n_83), .A1 (n_80), .A2 (n_81), .B1 (n_82), .B2 (M[27]));
INV_X1 i_110 (.ZN (n_82), .A (A[27]));
XNOR2_X1 i_109 (.ZN (p_0[27]), .A (n_80), .B (n_81));
XNOR2_X1 i_108 (.ZN (n_81), .A (A[27]), .B (M[27]));
OAI22_X1 i_107 (.ZN (n_80), .A1 (n_77), .A2 (n_78), .B1 (n_79), .B2 (A[26]));
INV_X1 i_106 (.ZN (n_79), .A (M[26]));
XNOR2_X1 i_105 (.ZN (p_0[26]), .A (n_77), .B (n_78));
XOR2_X1 i_104 (.Z (n_78), .A (A[26]), .B (M[26]));
AOI22_X1 i_103 (.ZN (n_77), .A1 (n_74), .A2 (n_75), .B1 (n_76), .B2 (M[25]));
INV_X1 i_102 (.ZN (n_76), .A (A[25]));
XNOR2_X1 i_101 (.ZN (p_0[25]), .A (n_74), .B (n_75));
XNOR2_X1 i_100 (.ZN (n_75), .A (A[25]), .B (M[25]));
OAI22_X1 i_99 (.ZN (n_74), .A1 (n_71), .A2 (n_72), .B1 (n_73), .B2 (A[24]));
INV_X1 i_98 (.ZN (n_73), .A (M[24]));
XNOR2_X1 i_97 (.ZN (p_0[24]), .A (n_71), .B (n_72));
XOR2_X1 i_96 (.Z (n_72), .A (A[24]), .B (M[24]));
AOI22_X1 i_95 (.ZN (n_71), .A1 (n_68), .A2 (n_69), .B1 (n_70), .B2 (M[23]));
INV_X1 i_94 (.ZN (n_70), .A (A[23]));
XNOR2_X1 i_93 (.ZN (p_0[23]), .A (n_68), .B (n_69));
XNOR2_X1 i_92 (.ZN (n_69), .A (A[23]), .B (M[23]));
OAI22_X1 i_91 (.ZN (n_68), .A1 (n_65), .A2 (n_66), .B1 (n_67), .B2 (A[22]));
INV_X1 i_90 (.ZN (n_67), .A (M[22]));
XNOR2_X1 i_89 (.ZN (p_0[22]), .A (n_65), .B (n_66));
XOR2_X1 i_88 (.Z (n_66), .A (A[22]), .B (M[22]));
AOI22_X1 i_87 (.ZN (n_65), .A1 (n_62), .A2 (n_63), .B1 (n_64), .B2 (M[21]));
INV_X1 i_86 (.ZN (n_64), .A (A[21]));
XNOR2_X1 i_85 (.ZN (p_0[21]), .A (n_62), .B (n_63));
XNOR2_X1 i_84 (.ZN (n_63), .A (A[21]), .B (M[21]));
OAI22_X1 i_83 (.ZN (n_62), .A1 (n_59), .A2 (n_60), .B1 (n_61), .B2 (A[20]));
INV_X1 i_82 (.ZN (n_61), .A (M[20]));
XNOR2_X1 i_81 (.ZN (p_0[20]), .A (n_59), .B (n_60));
XOR2_X1 i_80 (.Z (n_60), .A (A[20]), .B (M[20]));
AOI22_X1 i_79 (.ZN (n_59), .A1 (n_56), .A2 (n_57), .B1 (n_58), .B2 (M[19]));
INV_X1 i_78 (.ZN (n_58), .A (A[19]));
XNOR2_X1 i_77 (.ZN (p_0[19]), .A (n_56), .B (n_57));
XNOR2_X1 i_76 (.ZN (n_57), .A (A[19]), .B (M[19]));
OAI22_X1 i_75 (.ZN (n_56), .A1 (n_53), .A2 (n_54), .B1 (n_55), .B2 (A[18]));
INV_X1 i_74 (.ZN (n_55), .A (M[18]));
XNOR2_X1 i_73 (.ZN (p_0[18]), .A (n_53), .B (n_54));
XOR2_X1 i_72 (.Z (n_54), .A (A[18]), .B (M[18]));
AOI22_X1 i_71 (.ZN (n_53), .A1 (n_50), .A2 (n_51), .B1 (n_52), .B2 (M[17]));
INV_X1 i_70 (.ZN (n_52), .A (A[17]));
XNOR2_X1 i_69 (.ZN (p_0[17]), .A (n_50), .B (n_51));
XNOR2_X1 i_68 (.ZN (n_51), .A (A[17]), .B (M[17]));
OAI22_X1 i_67 (.ZN (n_50), .A1 (n_47), .A2 (n_48), .B1 (n_49), .B2 (A[16]));
INV_X1 i_66 (.ZN (n_49), .A (M[16]));
XNOR2_X1 i_65 (.ZN (p_0[16]), .A (n_47), .B (n_48));
XOR2_X1 i_64 (.Z (n_48), .A (A[16]), .B (M[16]));
AOI22_X1 i_63 (.ZN (n_47), .A1 (n_44), .A2 (n_45), .B1 (n_46), .B2 (M[15]));
INV_X1 i_62 (.ZN (n_46), .A (A[15]));
XNOR2_X1 i_61 (.ZN (p_0[15]), .A (n_44), .B (n_45));
XNOR2_X1 i_60 (.ZN (n_45), .A (A[15]), .B (M[15]));
OAI22_X1 i_59 (.ZN (n_44), .A1 (n_41), .A2 (n_42), .B1 (n_43), .B2 (A[14]));
INV_X1 i_58 (.ZN (n_43), .A (M[14]));
XNOR2_X1 i_57 (.ZN (p_0[14]), .A (n_41), .B (n_42));
XOR2_X1 i_56 (.Z (n_42), .A (A[14]), .B (M[14]));
AOI22_X1 i_55 (.ZN (n_41), .A1 (n_38), .A2 (n_39), .B1 (n_40), .B2 (M[13]));
INV_X1 i_54 (.ZN (n_40), .A (A[13]));
XNOR2_X1 i_53 (.ZN (p_0[13]), .A (n_38), .B (n_39));
XNOR2_X1 i_52 (.ZN (n_39), .A (A[13]), .B (M[13]));
OAI22_X1 i_51 (.ZN (n_38), .A1 (n_35), .A2 (n_36), .B1 (n_37), .B2 (A[12]));
INV_X1 i_50 (.ZN (n_37), .A (M[12]));
XNOR2_X1 i_49 (.ZN (p_0[12]), .A (n_35), .B (n_36));
XOR2_X1 i_48 (.Z (n_36), .A (A[12]), .B (M[12]));
AOI22_X1 i_47 (.ZN (n_35), .A1 (n_32), .A2 (n_33), .B1 (n_34), .B2 (M[11]));
INV_X1 i_46 (.ZN (n_34), .A (A[11]));
XNOR2_X1 i_45 (.ZN (p_0[11]), .A (n_32), .B (n_33));
XNOR2_X1 i_44 (.ZN (n_33), .A (A[11]), .B (M[11]));
OAI22_X1 i_43 (.ZN (n_32), .A1 (n_29), .A2 (n_30), .B1 (n_31), .B2 (A[10]));
INV_X1 i_42 (.ZN (n_31), .A (M[10]));
XNOR2_X1 i_41 (.ZN (p_0[10]), .A (n_29), .B (n_30));
XOR2_X1 i_40 (.Z (n_30), .A (A[10]), .B (M[10]));
AOI22_X1 i_39 (.ZN (n_29), .A1 (n_26), .A2 (n_27), .B1 (n_28), .B2 (M[9]));
INV_X1 i_38 (.ZN (n_28), .A (A[9]));
XNOR2_X1 i_37 (.ZN (p_0[9]), .A (n_26), .B (n_27));
XNOR2_X1 i_36 (.ZN (n_27), .A (A[9]), .B (M[9]));
OAI22_X1 i_35 (.ZN (n_26), .A1 (n_23), .A2 (n_24), .B1 (n_25), .B2 (A[8]));
INV_X1 i_34 (.ZN (n_25), .A (M[8]));
XNOR2_X1 i_33 (.ZN (p_0[8]), .A (n_23), .B (n_24));
XOR2_X1 i_32 (.Z (n_24), .A (A[8]), .B (M[8]));
AOI22_X1 i_31 (.ZN (n_23), .A1 (n_20), .A2 (n_21), .B1 (n_22), .B2 (M[7]));
INV_X1 i_30 (.ZN (n_22), .A (A[7]));
XNOR2_X1 i_29 (.ZN (p_0[7]), .A (n_20), .B (n_21));
XNOR2_X1 i_28 (.ZN (n_21), .A (A[7]), .B (M[7]));
OAI22_X1 i_27 (.ZN (n_20), .A1 (n_17), .A2 (n_18), .B1 (n_19), .B2 (A[6]));
INV_X1 i_26 (.ZN (n_19), .A (M[6]));
XNOR2_X1 i_25 (.ZN (p_0[6]), .A (n_17), .B (n_18));
XOR2_X1 i_24 (.Z (n_18), .A (A[6]), .B (M[6]));
AOI22_X1 i_23 (.ZN (n_17), .A1 (n_14), .A2 (n_15), .B1 (n_16), .B2 (M[5]));
INV_X1 i_22 (.ZN (n_16), .A (A[5]));
XNOR2_X1 i_21 (.ZN (p_0[5]), .A (n_14), .B (n_15));
XNOR2_X1 i_20 (.ZN (n_15), .A (A[5]), .B (M[5]));
OAI22_X1 i_19 (.ZN (n_14), .A1 (n_11), .A2 (n_12), .B1 (n_13), .B2 (A[4]));
INV_X1 i_18 (.ZN (n_13), .A (M[4]));
XNOR2_X1 i_17 (.ZN (p_0[4]), .A (n_11), .B (n_12));
XOR2_X1 i_16 (.Z (n_12), .A (A[4]), .B (M[4]));
AOI22_X1 i_15 (.ZN (n_11), .A1 (n_8), .A2 (n_9), .B1 (n_10), .B2 (M[3]));
INV_X1 i_14 (.ZN (n_10), .A (A[3]));
XNOR2_X1 i_13 (.ZN (p_0[3]), .A (n_8), .B (n_9));
XNOR2_X1 i_12 (.ZN (n_9), .A (A[3]), .B (M[3]));
OAI22_X1 i_11 (.ZN (n_8), .A1 (n_5), .A2 (n_6), .B1 (n_7), .B2 (A[2]));
INV_X1 i_10 (.ZN (n_7), .A (M[2]));
XNOR2_X1 i_9 (.ZN (p_0[2]), .A (n_5), .B (n_6));
XOR2_X1 i_8 (.Z (n_6), .A (M[2]), .B (A[2]));
AOI22_X1 i_7 (.ZN (n_5), .A1 (n_2), .A2 (n_3), .B1 (n_4), .B2 (M[1]));
INV_X1 i_6 (.ZN (n_4), .A (A[1]));
INV_X1 i_5 (.ZN (n_3), .A (n_1));
XOR2_X1 i_4 (.Z (p_0[1]), .A (n_2), .B (n_1));
XNOR2_X1 i_3 (.ZN (n_2), .A (A[1]), .B (M[1]));
OAI21_X1 i_2 (.ZN (p_0[0]), .A (n_1), .B1 (M[0]), .B2 (n_0));
NAND2_X1 i_1 (.ZN (n_1), .A1 (n_0), .A2 (M[0]));
INV_X1 i_0 (.ZN (n_0), .A (A[0]));

endmodule //datapath

module Booth (clk, rst, m, q, P);

output [63:0] P;
input clk;
input [31:0] m;
input [31:0] q;
input rst;
wire CTS_n178;
wire CLOCK_slh_n293;
wire CLOCK_slh_n373;
wire CLOCK_slh_n393;
wire CLOCK_slh_n383;
wire CLOCK_slh_n398;
wire CLOCK_slh_n368;
wire CLOCK_slh_n388;
wire CLOCK_slh_n378;
wire CLOCK_slh_n278;
wire CLOCK_slh_n273;
wire CLOCK_slh_n258;
wire CLOCK_slh_n253;
wire CLOCK_slh_n298;
wire CLOCK_slh_n248;
wire CLOCK_slh_n243;
wire CLOCK_slh_n268;
wire CLOCK_slh_n283;
wire CLOCK_slh_n333;
wire CLOCK_slh_n328;
wire CLOCK_slh_n263;
wire CLOCK_slh_n323;
wire CLOCK_slh_n318;
wire CLOCK_slh_n348;
wire CLOCK_slh_n303;
wire CLOCK_slh_n288;
wire CLOCK_slh_n343;
wire CLOCK_slh_n313;
wire CLOCK_slh_n338;
wire CLOCK_slh_n308;
wire CLOCK_slh_n353;
wire CLOCK_slh_n358;
wire CLOCK_slh_n363;
wire CTS_n105;
wire n_0_4;
wire n_0_5;
wire n_0_6;
wire n_0_7;
wire n_0_8;
wire n_0_9;
wire n_0_10;
wire n_0_11;
wire n_0_12;
wire n_0_13;
wire n_0_14;
wire n_0_15;
wire n_0_16;
wire n_0_17;
wire n_0_18;
wire n_0_19;
wire n_0_20;
wire n_0_21;
wire n_0_22;
wire n_0_23;
wire n_0_24;
wire n_0_25;
wire n_0_26;
wire n_0_27;
wire n_0_28;
wire n_0_29;
wire n_0_30;
wire n_0_31;
wire n_0_32;
wire n_0_33;
wire n_0_34;
wire n_0_35;
wire n_0_36;
wire n_0_37;
wire n_0_38;
wire n_0_39;
wire n_0_40;
wire n_0_41;
wire n_0_42;
wire n_0_43;
wire n_0_44;
wire n_0_45;
wire n_0_46;
wire n_0_47;
wire n_0_48;
wire n_0_49;
wire n_0_50;
wire n_0_51;
wire n_0_52;
wire n_0_53;
wire n_0_54;
wire n_0_55;
wire n_0_56;
wire n_0_57;
wire n_0_58;
wire n_0_59;
wire n_0_60;
wire n_0_61;
wire n_0_62;
wire n_0_63;
wire n_0_64;
wire n_0_65;
wire n_0_66;
wire n_0_67;
wire n_0_1;
wire n_0_0_0;
wire n_0_2;
wire n_0_0_1;
wire n_0_3;
wire n_0_0_2;
wire n_0_68;
wire n_0_0_3;
wire n_0_69;
wire n_0_0_4;
wire n_0_70;
wire n_0_0_5;
wire n_0_71;
wire n_0_0_6;
wire n_0_72;
wire n_0_0_7;
wire n_0_73;
wire n_0_0_8;
wire n_0_74;
wire n_0_0_9;
wire n_0_75;
wire n_0_0_10;
wire n_0_76;
wire n_0_0_11;
wire n_0_77;
wire n_0_0_12;
wire n_0_78;
wire n_0_0_13;
wire n_0_79;
wire n_0_0_14;
wire n_0_80;
wire n_0_0_15;
wire n_0_81;
wire n_0_0_16;
wire n_0_82;
wire n_0_0_17;
wire n_0_83;
wire n_0_0_18;
wire n_0_84;
wire n_0_0_19;
wire n_0_85;
wire n_0_0_20;
wire n_0_86;
wire n_0_0_21;
wire n_0_87;
wire n_0_0_22;
wire n_0_88;
wire n_0_0_23;
wire n_0_89;
wire n_0_0_24;
wire n_0_90;
wire n_0_0_25;
wire n_0_91;
wire n_0_0_26;
wire n_0_92;
wire n_0_0_27;
wire n_0_93;
wire n_0_0_28;
wire n_0_94;
wire n_0_0_29;
wire n_0_95;
wire n_0_0_30;
wire n_0_0_31;
wire n_0_114;
wire n_0_115;
wire n_0_116;
wire n_0_117;
wire n_0_118;
wire n_0_119;
wire n_0_120;
wire n_0_121;
wire n_0_122;
wire n_0_123;
wire n_0_124;
wire n_0_125;
wire n_0_126;
wire n_0_127;
wire n_0_128;
wire n_0_129;
wire n_0_130;
wire n_0_131;
wire n_0_132;
wire n_0_133;
wire n_0_134;
wire n_0_135;
wire n_0_136;
wire n_0_137;
wire n_0_138;
wire n_0_96;
wire n_0_97;
wire n_0_98;
wire n_0_99;
wire n_0_100;
wire n_0_101;
wire n_0_102;
wire n_0_0_32;
wire n_0_0_33;
wire n_0_0_34;
wire n_0_0_35;
wire n_0_0_36;
wire n_0_0_37;
wire n_0_107;
wire n_0_108;
wire n_0_0_38;
wire n_0_109;
wire n_0_0_39;
wire n_0_110;
wire n_0_0_40;
wire n_0_111;
wire n_0_0_41;
wire n_0_112;
wire n_0_0_42;
wire n_0_103;
wire n_0_104;
wire n_0_0_43;
wire n_0_0_44;
wire n_0_0_45;
wire n_0_0_46;
wire \Q[31] ;
wire \Q[30] ;
wire \Q[29] ;
wire \Q[28] ;
wire \Q[27] ;
wire \Q[26] ;
wire \Q[25] ;
wire \Q[24] ;
wire \Q[23] ;
wire \Q[22] ;
wire \Q[21] ;
wire \Q[20] ;
wire \Q[19] ;
wire \Q[18] ;
wire \Q[17] ;
wire \Q[16] ;
wire \Q[15] ;
wire \Q[14] ;
wire \Q[13] ;
wire \Q[12] ;
wire \Q[11] ;
wire \Q[10] ;
wire \Q[9] ;
wire \Q[8] ;
wire \Q[7] ;
wire \Q[6] ;
wire \Q[5] ;
wire \Q[4] ;
wire \Q[3] ;
wire \Q[2] ;
wire \Q[1] ;
wire \Q[0] ;
wire \A[31] ;
wire \A[29] ;
wire \A[28] ;
wire \A[27] ;
wire \A[26] ;
wire \A[25] ;
wire \A[24] ;
wire \A[23] ;
wire \A[22] ;
wire \A[21] ;
wire \A[20] ;
wire \A[19] ;
wire \A[18] ;
wire \A[17] ;
wire \A[16] ;
wire \A[15] ;
wire \A[14] ;
wire \A[13] ;
wire \A[12] ;
wire \A[11] ;
wire \A[10] ;
wire \A[9] ;
wire \A[8] ;
wire \A[7] ;
wire \A[6] ;
wire \A[5] ;
wire \A[4] ;
wire \A[3] ;
wire \A[2] ;
wire \A[1] ;
wire \A[0] ;
wire CTS_n106;
wire \M[31] ;
wire \M[30] ;
wire \M[29] ;
wire \M[28] ;
wire \M[27] ;
wire \M[26] ;
wire \M[25] ;
wire \M[24] ;
wire \M[23] ;
wire \M[22] ;
wire \M[21] ;
wire \M[20] ;
wire \M[19] ;
wire \M[18] ;
wire \M[17] ;
wire \M[16] ;
wire \M[15] ;
wire \M[14] ;
wire \M[13] ;
wire \M[12] ;
wire \M[11] ;
wire \M[10] ;
wire \M[9] ;
wire \M[8] ;
wire \M[7] ;
wire \M[6] ;
wire \M[5] ;
wire \M[4] ;
wire \M[3] ;
wire \M[2] ;
wire \M[1] ;
wire \M[0] ;
wire q1;
wire \n[5] ;
wire \n[4] ;
wire \n[3] ;
wire \n[2] ;
wire \n[1] ;
wire \n[0] ;
wire CTS_n8;
wire n_0_113;
wire uc_0;
wire uc_1;
wire drc_ipo_n6;
wire drc_ipo_n5;
wire CTS_n9;
wire CTS_n214;
wire CTS_n101;
wire CTS_n56;
wire CTS_n193;

// WARNING . Detected multiport output net(s). Introducing ASSIGN statements.
// This may cause simulation/synthesis mismatches . 
assign P[63] = P[62];

INV_X1 i_0_12 (.ZN (n_0_113), .A (n_0_104));
CLKGATETST_X8 clk_gate_A_reg (.GCK (CTS_n56), .CK (CTS_n193), .E (n_0_113), .SE (1'b0 ));
DFF_X1 \n_reg[0]  (.Q (\n[0] ), .CK (CTS_n8), .D (n_0_107));
DFF_X1 \n_reg[1]  (.Q (\n[1] ), .CK (CTS_n8), .D (n_0_108));
DFF_X1 \n_reg[2]  (.Q (\n[2] ), .CK (CTS_n8), .D (n_0_109));
DFF_X1 \n_reg[3]  (.Q (\n[3] ), .CK (CTS_n8), .D (n_0_110));
DFF_X1 \n_reg[4]  (.Q (\n[4] ), .CK (CTS_n8), .D (n_0_111));
DFF_X1 \n_reg[5]  (.Q (\n[5] ), .CK (CTS_n8), .D (n_0_112));
DFF_X1 q1_reg (.Q (q1), .CK (CTS_n8), .D (n_0_103));
DFF_X1 \M_reg[0]  (.Q (\M[0] ), .CK (CTS_n101), .D (CLOCK_slh_n363));
DFF_X1 \M_reg[1]  (.Q (\M[1] ), .CK (CTS_n101), .D (CLOCK_slh_n358));
DFF_X1 \M_reg[2]  (.Q (\M[2] ), .CK (CTS_n101), .D (CLOCK_slh_n353));
DFF_X1 \M_reg[3]  (.Q (\M[3] ), .CK (CTS_n101), .D (CLOCK_slh_n308));
DFF_X1 \M_reg[4]  (.Q (\M[4] ), .CK (CTS_n101), .D (CLOCK_slh_n338));
DFF_X1 \M_reg[5]  (.Q (\M[5] ), .CK (CTS_n101), .D (CLOCK_slh_n313));
DFF_X1 \M_reg[6]  (.Q (\M[6] ), .CK (CTS_n101), .D (CLOCK_slh_n343));
DFF_X1 \M_reg[7]  (.Q (\M[7] ), .CK (CTS_n101), .D (CLOCK_slh_n288));
DFF_X1 \M_reg[8]  (.Q (\M[8] ), .CK (CTS_n101), .D (CLOCK_slh_n303));
DFF_X1 \M_reg[9]  (.Q (\M[9] ), .CK (CTS_n101), .D (CLOCK_slh_n348));
DFF_X1 \M_reg[10]  (.Q (\M[10] ), .CK (CTS_n101), .D (CLOCK_slh_n318));
DFF_X1 \M_reg[11]  (.Q (\M[11] ), .CK (CTS_n101), .D (CLOCK_slh_n323));
DFF_X1 \M_reg[12]  (.Q (\M[12] ), .CK (CTS_n101), .D (CLOCK_slh_n263));
DFF_X1 \M_reg[13]  (.Q (\M[13] ), .CK (CTS_n101), .D (CLOCK_slh_n328));
DFF_X1 \M_reg[14]  (.Q (\M[14] ), .CK (CTS_n101), .D (CLOCK_slh_n333));
DFF_X1 \M_reg[15]  (.Q (\M[15] ), .CK (CTS_n101), .D (CLOCK_slh_n283));
DFF_X1 \M_reg[16]  (.Q (\M[16] ), .CK (CTS_n101), .D (CLOCK_slh_n268));
DFF_X1 \M_reg[17]  (.Q (\M[17] ), .CK (CTS_n101), .D (CLOCK_slh_n243));
DFF_X1 \M_reg[18]  (.Q (\M[18] ), .CK (CTS_n101), .D (CLOCK_slh_n248));
DFF_X1 \M_reg[19]  (.Q (\M[19] ), .CK (CTS_n101), .D (CLOCK_slh_n298));
DFF_X1 \M_reg[20]  (.Q (\M[20] ), .CK (CTS_n101), .D (CLOCK_slh_n253));
DFF_X1 \M_reg[21]  (.Q (\M[21] ), .CK (CTS_n101), .D (CLOCK_slh_n258));
DFF_X1 \M_reg[22]  (.Q (\M[22] ), .CK (CTS_n101), .D (CLOCK_slh_n273));
DFF_X1 \M_reg[23]  (.Q (\M[23] ), .CK (CTS_n101), .D (CLOCK_slh_n278));
DFF_X1 \M_reg[24]  (.Q (\M[24] ), .CK (CTS_n101), .D (CLOCK_slh_n378));
DFF_X1 \M_reg[25]  (.Q (\M[25] ), .CK (CTS_n101), .D (CLOCK_slh_n388));
DFF_X1 \M_reg[26]  (.Q (\M[26] ), .CK (CTS_n101), .D (CLOCK_slh_n368));
DFF_X1 \M_reg[27]  (.Q (\M[27] ), .CK (CTS_n101), .D (CLOCK_slh_n398));
DFF_X1 \M_reg[28]  (.Q (\M[28] ), .CK (CTS_n101), .D (CLOCK_slh_n383));
DFF_X1 \M_reg[29]  (.Q (\M[29] ), .CK (CTS_n101), .D (CLOCK_slh_n393));
DFF_X1 \M_reg[30]  (.Q (\M[30] ), .CK (CTS_n101), .D (CLOCK_slh_n373));
DFF_X1 \M_reg[31]  (.Q (\M[31] ), .CK (CTS_n101), .D (CLOCK_slh_n293));
CLKGATETST_X8 clk_gate_M_reg (.GCK (CTS_n101), .CK (CTS_n178), .E (rst), .SE (1'b0 ));
DFF_X1 \A_reg[0]  (.Q (\A[0] ), .CK (CTS_n8), .D (n_0_1));
DFF_X1 \A_reg[1]  (.Q (\A[1] ), .CK (CTS_n8), .D (n_0_2));
DFF_X1 \A_reg[2]  (.Q (\A[2] ), .CK (CTS_n8), .D (n_0_3));
DFF_X1 \A_reg[3]  (.Q (\A[3] ), .CK (CTS_n8), .D (n_0_68));
DFF_X1 \A_reg[4]  (.Q (\A[4] ), .CK (CTS_n9), .D (n_0_69));
DFF_X1 \A_reg[5]  (.Q (\A[5] ), .CK (CTS_n9), .D (n_0_70));
DFF_X1 \A_reg[6]  (.Q (\A[6] ), .CK (CTS_n9), .D (n_0_71));
DFF_X1 \A_reg[7]  (.Q (\A[7] ), .CK (CTS_n9), .D (n_0_72));
DFF_X1 \A_reg[8]  (.Q (\A[8] ), .CK (CTS_n9), .D (n_0_73));
DFF_X1 \A_reg[9]  (.Q (\A[9] ), .CK (CTS_n9), .D (n_0_74));
DFF_X1 \A_reg[10]  (.Q (\A[10] ), .CK (CTS_n9), .D (n_0_75));
DFF_X1 \A_reg[11]  (.Q (\A[11] ), .CK (CTS_n9), .D (n_0_76));
DFF_X1 \A_reg[12]  (.Q (\A[12] ), .CK (CTS_n9), .D (n_0_77));
DFF_X1 \A_reg[13]  (.Q (\A[13] ), .CK (CTS_n9), .D (n_0_78));
DFF_X1 \A_reg[14]  (.Q (\A[14] ), .CK (CTS_n9), .D (n_0_79));
DFF_X1 \A_reg[15]  (.Q (\A[15] ), .CK (CTS_n9), .D (n_0_80));
DFF_X1 \A_reg[16]  (.Q (\A[16] ), .CK (CTS_n9), .D (n_0_81));
DFF_X1 \A_reg[17]  (.Q (\A[17] ), .CK (CTS_n9), .D (n_0_82));
DFF_X1 \A_reg[18]  (.Q (\A[18] ), .CK (CTS_n9), .D (n_0_83));
DFF_X1 \A_reg[19]  (.Q (\A[19] ), .CK (CTS_n9), .D (n_0_84));
DFF_X1 \A_reg[20]  (.Q (\A[20] ), .CK (CTS_n9), .D (n_0_85));
DFF_X1 \A_reg[21]  (.Q (\A[21] ), .CK (CTS_n9), .D (n_0_86));
DFF_X1 \A_reg[22]  (.Q (\A[22] ), .CK (CTS_n9), .D (n_0_87));
DFF_X1 \A_reg[23]  (.Q (\A[23] ), .CK (CTS_n9), .D (n_0_88));
DFF_X1 \A_reg[24]  (.Q (\A[24] ), .CK (CTS_n9), .D (n_0_89));
DFF_X1 \A_reg[25]  (.Q (\A[25] ), .CK (CTS_n8), .D (n_0_90));
DFF_X1 \A_reg[26]  (.Q (\A[26] ), .CK (CTS_n8), .D (n_0_91));
DFF_X1 \A_reg[27]  (.Q (\A[27] ), .CK (CTS_n8), .D (n_0_92));
DFF_X1 \A_reg[28]  (.Q (\A[28] ), .CK (CTS_n8), .D (n_0_93));
DFF_X1 \A_reg[29]  (.Q (\A[29] ), .CK (CTS_n8), .D (n_0_94));
DFF_X1 \A_reg[31]  (.Q (\A[31] ), .CK (CTS_n8), .D (n_0_95));
DFF_X1 \Q_reg[0]  (.Q (\Q[0] ), .CK (CTS_n8), .D (n_0_114));
DFF_X1 \Q_reg[1]  (.Q (\Q[1] ), .CK (CTS_n8), .D (n_0_115));
DFF_X1 \Q_reg[2]  (.Q (\Q[2] ), .CK (CTS_n8), .D (n_0_116));
DFF_X1 \Q_reg[3]  (.Q (\Q[3] ), .CK (CTS_n9), .D (n_0_117));
DFF_X1 \Q_reg[4]  (.Q (\Q[4] ), .CK (CTS_n9), .D (n_0_118));
DFF_X1 \Q_reg[5]  (.Q (\Q[5] ), .CK (CTS_n9), .D (n_0_119));
DFF_X1 \Q_reg[6]  (.Q (\Q[6] ), .CK (CTS_n9), .D (n_0_120));
DFF_X1 \Q_reg[7]  (.Q (\Q[7] ), .CK (CTS_n9), .D (n_0_121));
DFF_X1 \Q_reg[8]  (.Q (\Q[8] ), .CK (CTS_n9), .D (n_0_122));
DFF_X1 \Q_reg[9]  (.Q (\Q[9] ), .CK (CTS_n9), .D (n_0_123));
DFF_X1 \Q_reg[10]  (.Q (\Q[10] ), .CK (CTS_n9), .D (n_0_124));
DFF_X1 \Q_reg[11]  (.Q (\Q[11] ), .CK (CTS_n9), .D (n_0_125));
DFF_X1 \Q_reg[12]  (.Q (\Q[12] ), .CK (CTS_n9), .D (n_0_126));
DFF_X1 \Q_reg[13]  (.Q (\Q[13] ), .CK (CTS_n9), .D (n_0_127));
DFF_X1 \Q_reg[14]  (.Q (\Q[14] ), .CK (CTS_n9), .D (n_0_128));
DFF_X1 \Q_reg[15]  (.Q (\Q[15] ), .CK (CTS_n8), .D (n_0_129));
DFF_X1 \Q_reg[16]  (.Q (\Q[16] ), .CK (CTS_n8), .D (n_0_130));
DFF_X1 \Q_reg[17]  (.Q (\Q[17] ), .CK (CTS_n8), .D (n_0_131));
DFF_X1 \Q_reg[18]  (.Q (\Q[18] ), .CK (CTS_n8), .D (n_0_132));
DFF_X1 \Q_reg[19]  (.Q (\Q[19] ), .CK (CTS_n8), .D (n_0_133));
DFF_X1 \Q_reg[20]  (.Q (\Q[20] ), .CK (CTS_n8), .D (n_0_134));
DFF_X1 \Q_reg[21]  (.Q (\Q[21] ), .CK (CTS_n8), .D (n_0_135));
DFF_X1 \Q_reg[22]  (.Q (\Q[22] ), .CK (CTS_n8), .D (n_0_136));
DFF_X1 \Q_reg[23]  (.Q (\Q[23] ), .CK (CTS_n8), .D (n_0_137));
DFF_X1 \Q_reg[24]  (.Q (\Q[24] ), .CK (CTS_n8), .D (n_0_138));
DFF_X1 \Q_reg[25]  (.Q (\Q[25] ), .CK (CTS_n8), .D (n_0_96));
DFF_X1 \Q_reg[26]  (.Q (\Q[26] ), .CK (CTS_n8), .D (n_0_97));
DFF_X1 \Q_reg[27]  (.Q (\Q[27] ), .CK (CTS_n8), .D (n_0_98));
DFF_X1 \Q_reg[28]  (.Q (\Q[28] ), .CK (CTS_n8), .D (n_0_99));
DFF_X1 \Q_reg[29]  (.Q (\Q[29] ), .CK (CTS_n8), .D (n_0_100));
DFF_X1 \Q_reg[30]  (.Q (\Q[30] ), .CK (CTS_n8), .D (n_0_101));
DFF_X1 \Q_reg[31]  (.Q (\Q[31] ), .CK (CTS_n8), .D (n_0_102));
INV_X1 i_0_0_117 (.ZN (n_0_0_46), .A (q1));
INV_X1 i_0_0_116 (.ZN (n_0_0_45), .A (\Q[0] ));
OR3_X1 i_0_0_115 (.ZN (n_0_0_44), .A1 (\n[2] ), .A2 (\n[1] ), .A3 (\n[0] ));
OR3_X1 i_0_0_114 (.ZN (n_0_0_43), .A1 (n_0_0_44), .A2 (\n[3] ), .A3 (\n[4] ));
NOR3_X1 i_0_0_113 (.ZN (n_0_104), .A1 (n_0_0_43), .A2 (rst), .A3 (\n[5] ));
NOR2_X1 i_0_0_112 (.ZN (n_0_103), .A1 (n_0_0_45), .A2 (rst));
AOI21_X1 i_0_0_111 (.ZN (n_0_0_42), .A (rst), .B1 (n_0_0_43), .B2 (\n[5] ));
OAI21_X1 i_0_0_110 (.ZN (n_0_112), .A (n_0_0_42), .B1 (n_0_0_43), .B2 (\n[5] ));
OAI21_X1 i_0_0_109 (.ZN (n_0_0_41), .A (\n[4] ), .B1 (n_0_0_44), .B2 (\n[3] ));
AOI21_X1 i_0_0_108 (.ZN (n_0_111), .A (rst), .B1 (n_0_0_43), .B2 (n_0_0_41));
XOR2_X1 i_0_0_107 (.Z (n_0_0_40), .A (\n[3] ), .B (n_0_0_44));
NOR2_X1 i_0_0_106 (.ZN (n_0_110), .A1 (rst), .A2 (n_0_0_40));
OAI21_X1 i_0_0_105 (.ZN (n_0_0_39), .A (\n[2] ), .B1 (\n[1] ), .B2 (\n[0] ));
AOI21_X1 i_0_0_104 (.ZN (n_0_109), .A (rst), .B1 (n_0_0_44), .B2 (n_0_0_39));
XOR2_X1 i_0_0_103 (.Z (n_0_0_38), .A (\n[1] ), .B (\n[0] ));
NOR2_X1 i_0_0_102 (.ZN (n_0_108), .A1 (rst), .A2 (n_0_0_38));
NOR2_X1 i_0_0_101 (.ZN (n_0_107), .A1 (\n[0] ), .A2 (rst));
XNOR2_X1 i_0_0_100 (.ZN (n_0_0_37), .A (n_0_0_46), .B (\Q[0] ));
NOR2_X4 i_0_0_99 (.ZN (n_0_0_36), .A1 (n_0_0_37), .A2 (rst));
NAND2_X1 i_0_0_98 (.ZN (n_0_0_35), .A1 (\A[0] ), .A2 (n_0_0_36));
NOR3_X1 i_0_0_97 (.ZN (n_0_0_34), .A1 (n_0_0_46), .A2 (\Q[0] ), .A3 (rst));
NOR3_X1 i_0_0_96 (.ZN (n_0_0_33), .A1 (n_0_0_45), .A2 (q1), .A3 (rst));
AOI222_X1 i_0_0_95 (.ZN (n_0_0_32), .A1 (rst), .A2 (q[31]), .B1 (drc_ipo_n5), .B2 (n_0_36)
    , .C1 (drc_ipo_n6), .C2 (n_0_4));
NAND2_X1 i_0_0_94 (.ZN (n_0_102), .A1 (n_0_0_32), .A2 (n_0_0_35));
MUX2_X1 i_0_0_93 (.Z (n_0_101), .A (\Q[31] ), .B (q[30]), .S (rst));
MUX2_X1 i_0_0_92 (.Z (n_0_100), .A (\Q[30] ), .B (q[29]), .S (rst));
MUX2_X1 i_0_0_91 (.Z (n_0_99), .A (\Q[29] ), .B (q[28]), .S (rst));
MUX2_X1 i_0_0_90 (.Z (n_0_98), .A (\Q[28] ), .B (q[27]), .S (rst));
MUX2_X1 i_0_0_89 (.Z (n_0_97), .A (\Q[27] ), .B (q[26]), .S (rst));
MUX2_X1 i_0_0_88 (.Z (n_0_96), .A (\Q[26] ), .B (q[25]), .S (rst));
MUX2_X1 i_0_0_87 (.Z (n_0_138), .A (\Q[25] ), .B (q[24]), .S (rst));
MUX2_X1 i_0_0_86 (.Z (n_0_137), .A (\Q[24] ), .B (q[23]), .S (rst));
MUX2_X1 i_0_0_85 (.Z (n_0_136), .A (\Q[23] ), .B (q[22]), .S (rst));
MUX2_X1 i_0_0_84 (.Z (n_0_135), .A (\Q[22] ), .B (q[21]), .S (rst));
MUX2_X1 i_0_0_83 (.Z (n_0_134), .A (\Q[21] ), .B (q[20]), .S (rst));
MUX2_X1 i_0_0_82 (.Z (n_0_133), .A (\Q[20] ), .B (q[19]), .S (rst));
MUX2_X1 i_0_0_81 (.Z (n_0_132), .A (\Q[19] ), .B (q[18]), .S (rst));
MUX2_X1 i_0_0_80 (.Z (n_0_131), .A (\Q[18] ), .B (q[17]), .S (rst));
MUX2_X1 i_0_0_79 (.Z (n_0_130), .A (\Q[17] ), .B (q[16]), .S (rst));
MUX2_X1 i_0_0_78 (.Z (n_0_129), .A (\Q[16] ), .B (q[15]), .S (rst));
MUX2_X1 i_0_0_77 (.Z (n_0_128), .A (\Q[15] ), .B (q[14]), .S (rst));
MUX2_X1 i_0_0_76 (.Z (n_0_127), .A (\Q[14] ), .B (q[13]), .S (rst));
MUX2_X1 i_0_0_75 (.Z (n_0_126), .A (\Q[13] ), .B (q[12]), .S (rst));
MUX2_X1 i_0_0_74 (.Z (n_0_125), .A (\Q[12] ), .B (q[11]), .S (rst));
MUX2_X1 i_0_0_73 (.Z (n_0_124), .A (\Q[11] ), .B (q[10]), .S (rst));
MUX2_X1 i_0_0_72 (.Z (n_0_123), .A (\Q[10] ), .B (q[9]), .S (rst));
MUX2_X1 i_0_0_71 (.Z (n_0_122), .A (\Q[9] ), .B (q[8]), .S (rst));
MUX2_X1 i_0_0_70 (.Z (n_0_121), .A (\Q[8] ), .B (q[7]), .S (rst));
MUX2_X1 i_0_0_69 (.Z (n_0_120), .A (\Q[7] ), .B (q[6]), .S (rst));
MUX2_X1 i_0_0_68 (.Z (n_0_119), .A (\Q[6] ), .B (q[5]), .S (rst));
MUX2_X1 i_0_0_67 (.Z (n_0_118), .A (\Q[5] ), .B (q[4]), .S (rst));
MUX2_X1 i_0_0_66 (.Z (n_0_117), .A (\Q[4] ), .B (q[3]), .S (rst));
MUX2_X1 i_0_0_65 (.Z (n_0_116), .A (\Q[3] ), .B (q[2]), .S (rst));
MUX2_X1 i_0_0_64 (.Z (n_0_115), .A (\Q[2] ), .B (q[1]), .S (rst));
MUX2_X1 i_0_0_63 (.Z (n_0_114), .A (\Q[1] ), .B (q[0]), .S (rst));
NAND2_X1 i_0_0_62 (.ZN (n_0_0_31), .A1 (\A[31] ), .A2 (n_0_0_36));
AOI22_X1 i_0_0_61 (.ZN (n_0_0_30), .A1 (n_0_67), .A2 (drc_ipo_n5), .B1 (drc_ipo_n6), .B2 (n_0_35));
NAND2_X1 i_0_0_60 (.ZN (n_0_95), .A1 (n_0_0_31), .A2 (n_0_0_30));
AOI22_X1 i_0_0_59 (.ZN (n_0_0_29), .A1 (n_0_66), .A2 (drc_ipo_n5), .B1 (drc_ipo_n6), .B2 (n_0_34));
NAND2_X1 i_0_0_58 (.ZN (n_0_94), .A1 (n_0_0_31), .A2 (n_0_0_29));
AOI222_X1 i_0_0_57 (.ZN (n_0_0_28), .A1 (\A[29] ), .A2 (n_0_0_36), .B1 (drc_ipo_n5)
    , .B2 (n_0_65), .C1 (drc_ipo_n6), .C2 (n_0_33));
INV_X1 i_0_0_56 (.ZN (n_0_93), .A (n_0_0_28));
AOI222_X1 i_0_0_55 (.ZN (n_0_0_27), .A1 (\A[28] ), .A2 (n_0_0_36), .B1 (drc_ipo_n5)
    , .B2 (n_0_64), .C1 (drc_ipo_n6), .C2 (n_0_32));
INV_X1 i_0_0_54 (.ZN (n_0_92), .A (n_0_0_27));
AOI222_X1 i_0_0_53 (.ZN (n_0_0_26), .A1 (\A[27] ), .A2 (n_0_0_36), .B1 (drc_ipo_n5)
    , .B2 (n_0_63), .C1 (drc_ipo_n6), .C2 (n_0_31));
INV_X1 i_0_0_52 (.ZN (n_0_91), .A (n_0_0_26));
AOI222_X1 i_0_0_51 (.ZN (n_0_0_25), .A1 (\A[26] ), .A2 (n_0_0_36), .B1 (drc_ipo_n5)
    , .B2 (n_0_62), .C1 (drc_ipo_n6), .C2 (n_0_30));
INV_X1 i_0_0_50 (.ZN (n_0_90), .A (n_0_0_25));
AOI222_X1 i_0_0_49 (.ZN (n_0_0_24), .A1 (\A[25] ), .A2 (n_0_0_36), .B1 (drc_ipo_n5)
    , .B2 (n_0_61), .C1 (drc_ipo_n6), .C2 (n_0_29));
INV_X1 i_0_0_48 (.ZN (n_0_89), .A (n_0_0_24));
AOI222_X1 i_0_0_47 (.ZN (n_0_0_23), .A1 (\A[24] ), .A2 (n_0_0_36), .B1 (drc_ipo_n5)
    , .B2 (n_0_60), .C1 (drc_ipo_n6), .C2 (n_0_28));
INV_X1 i_0_0_46 (.ZN (n_0_88), .A (n_0_0_23));
AOI222_X1 i_0_0_45 (.ZN (n_0_0_22), .A1 (\A[23] ), .A2 (n_0_0_36), .B1 (drc_ipo_n5)
    , .B2 (n_0_59), .C1 (drc_ipo_n6), .C2 (n_0_27));
INV_X1 i_0_0_44 (.ZN (n_0_87), .A (n_0_0_22));
AOI222_X1 i_0_0_43 (.ZN (n_0_0_21), .A1 (\A[22] ), .A2 (n_0_0_36), .B1 (drc_ipo_n5)
    , .B2 (n_0_58), .C1 (drc_ipo_n6), .C2 (n_0_26));
INV_X1 i_0_0_42 (.ZN (n_0_86), .A (n_0_0_21));
AOI222_X1 i_0_0_41 (.ZN (n_0_0_20), .A1 (\A[21] ), .A2 (n_0_0_36), .B1 (drc_ipo_n5)
    , .B2 (n_0_57), .C1 (drc_ipo_n6), .C2 (n_0_25));
INV_X1 i_0_0_40 (.ZN (n_0_85), .A (n_0_0_20));
AOI222_X1 i_0_0_39 (.ZN (n_0_0_19), .A1 (\A[20] ), .A2 (n_0_0_36), .B1 (drc_ipo_n5)
    , .B2 (n_0_56), .C1 (drc_ipo_n6), .C2 (n_0_24));
INV_X1 i_0_0_38 (.ZN (n_0_84), .A (n_0_0_19));
AOI222_X1 i_0_0_37 (.ZN (n_0_0_18), .A1 (\A[19] ), .A2 (n_0_0_36), .B1 (drc_ipo_n5)
    , .B2 (n_0_55), .C1 (drc_ipo_n6), .C2 (n_0_23));
INV_X1 i_0_0_36 (.ZN (n_0_83), .A (n_0_0_18));
AOI222_X1 i_0_0_35 (.ZN (n_0_0_17), .A1 (\A[18] ), .A2 (n_0_0_36), .B1 (drc_ipo_n5)
    , .B2 (n_0_54), .C1 (drc_ipo_n6), .C2 (n_0_22));
INV_X1 i_0_0_34 (.ZN (n_0_82), .A (n_0_0_17));
AOI222_X1 i_0_0_33 (.ZN (n_0_0_16), .A1 (\A[17] ), .A2 (n_0_0_36), .B1 (drc_ipo_n5)
    , .B2 (n_0_53), .C1 (drc_ipo_n6), .C2 (n_0_21));
INV_X1 i_0_0_32 (.ZN (n_0_81), .A (n_0_0_16));
AOI222_X1 i_0_0_31 (.ZN (n_0_0_15), .A1 (\A[16] ), .A2 (n_0_0_36), .B1 (drc_ipo_n5)
    , .B2 (n_0_52), .C1 (drc_ipo_n6), .C2 (n_0_20));
INV_X1 i_0_0_30 (.ZN (n_0_80), .A (n_0_0_15));
AOI222_X1 i_0_0_29 (.ZN (n_0_0_14), .A1 (\A[15] ), .A2 (n_0_0_36), .B1 (drc_ipo_n5)
    , .B2 (n_0_51), .C1 (drc_ipo_n6), .C2 (n_0_19));
INV_X1 i_0_0_28 (.ZN (n_0_79), .A (n_0_0_14));
AOI222_X1 i_0_0_27 (.ZN (n_0_0_13), .A1 (\A[14] ), .A2 (n_0_0_36), .B1 (drc_ipo_n5)
    , .B2 (n_0_50), .C1 (drc_ipo_n6), .C2 (n_0_18));
INV_X1 i_0_0_26 (.ZN (n_0_78), .A (n_0_0_13));
AOI222_X1 i_0_0_25 (.ZN (n_0_0_12), .A1 (\A[13] ), .A2 (n_0_0_36), .B1 (drc_ipo_n5)
    , .B2 (n_0_49), .C1 (drc_ipo_n6), .C2 (n_0_17));
INV_X1 i_0_0_24 (.ZN (n_0_77), .A (n_0_0_12));
AOI222_X1 i_0_0_23 (.ZN (n_0_0_11), .A1 (\A[12] ), .A2 (n_0_0_36), .B1 (drc_ipo_n5)
    , .B2 (n_0_48), .C1 (drc_ipo_n6), .C2 (n_0_16));
INV_X1 i_0_0_22 (.ZN (n_0_76), .A (n_0_0_11));
AOI222_X1 i_0_0_21 (.ZN (n_0_0_10), .A1 (\A[11] ), .A2 (n_0_0_36), .B1 (drc_ipo_n5)
    , .B2 (n_0_47), .C1 (drc_ipo_n6), .C2 (n_0_15));
INV_X1 i_0_0_20 (.ZN (n_0_75), .A (n_0_0_10));
AOI222_X1 i_0_0_19 (.ZN (n_0_0_9), .A1 (\A[10] ), .A2 (n_0_0_36), .B1 (drc_ipo_n5)
    , .B2 (n_0_46), .C1 (drc_ipo_n6), .C2 (n_0_14));
INV_X1 i_0_0_18 (.ZN (n_0_74), .A (n_0_0_9));
AOI222_X1 i_0_0_17 (.ZN (n_0_0_8), .A1 (\A[9] ), .A2 (n_0_0_36), .B1 (drc_ipo_n5)
    , .B2 (n_0_45), .C1 (drc_ipo_n6), .C2 (n_0_13));
INV_X1 i_0_0_16 (.ZN (n_0_73), .A (n_0_0_8));
AOI222_X1 i_0_0_15 (.ZN (n_0_0_7), .A1 (\A[8] ), .A2 (n_0_0_36), .B1 (drc_ipo_n5)
    , .B2 (n_0_44), .C1 (drc_ipo_n6), .C2 (n_0_12));
INV_X1 i_0_0_14 (.ZN (n_0_72), .A (n_0_0_7));
AOI222_X1 i_0_0_13 (.ZN (n_0_0_6), .A1 (\A[7] ), .A2 (n_0_0_36), .B1 (drc_ipo_n5)
    , .B2 (n_0_43), .C1 (drc_ipo_n6), .C2 (n_0_11));
INV_X1 i_0_0_12 (.ZN (n_0_71), .A (n_0_0_6));
AOI222_X1 i_0_0_11 (.ZN (n_0_0_5), .A1 (\A[6] ), .A2 (n_0_0_36), .B1 (drc_ipo_n5)
    , .B2 (n_0_42), .C1 (drc_ipo_n6), .C2 (n_0_10));
INV_X1 i_0_0_10 (.ZN (n_0_70), .A (n_0_0_5));
AOI222_X1 i_0_0_9 (.ZN (n_0_0_4), .A1 (\A[5] ), .A2 (n_0_0_36), .B1 (drc_ipo_n5), .B2 (n_0_41)
    , .C1 (drc_ipo_n6), .C2 (n_0_9));
INV_X1 i_0_0_8 (.ZN (n_0_69), .A (n_0_0_4));
AOI222_X1 i_0_0_7 (.ZN (n_0_0_3), .A1 (\A[4] ), .A2 (n_0_0_36), .B1 (drc_ipo_n5), .B2 (n_0_40)
    , .C1 (drc_ipo_n6), .C2 (n_0_8));
INV_X1 i_0_0_6 (.ZN (n_0_68), .A (n_0_0_3));
AOI222_X1 i_0_0_5 (.ZN (n_0_0_2), .A1 (\A[3] ), .A2 (n_0_0_36), .B1 (drc_ipo_n5), .B2 (n_0_39)
    , .C1 (drc_ipo_n6), .C2 (n_0_7));
INV_X1 i_0_0_4 (.ZN (n_0_3), .A (n_0_0_2));
AOI222_X1 i_0_0_3 (.ZN (n_0_0_1), .A1 (\A[2] ), .A2 (n_0_0_36), .B1 (drc_ipo_n5), .B2 (n_0_38)
    , .C1 (drc_ipo_n6), .C2 (n_0_6));
INV_X1 i_0_0_2 (.ZN (n_0_2), .A (n_0_0_1));
AOI222_X1 i_0_0_1 (.ZN (n_0_0_0), .A1 (\A[1] ), .A2 (n_0_0_36), .B1 (drc_ipo_n5), .B2 (n_0_37)
    , .C1 (drc_ipo_n6), .C2 (n_0_5));
INV_X1 i_0_0_0 (.ZN (n_0_1), .A (n_0_0_0));
datapath__0_1 i_0_4 (.p_0 ({n_0_67, n_0_66, n_0_65, n_0_64, n_0_63, n_0_62, n_0_61, 
    n_0_60, n_0_59, n_0_58, n_0_57, n_0_56, n_0_55, n_0_54, n_0_53, n_0_52, n_0_51, 
    n_0_50, n_0_49, n_0_48, n_0_47, n_0_46, n_0_45, n_0_44, n_0_43, n_0_42, n_0_41, 
    n_0_40, n_0_39, n_0_38, n_0_37, n_0_36}), .A ({\A[31] , uc_1, \A[29] , \A[28] , 
    \A[27] , \A[26] , \A[25] , \A[24] , \A[23] , \A[22] , \A[21] , \A[20] , \A[19] , 
    \A[18] , \A[17] , \A[16] , \A[15] , \A[14] , \A[13] , \A[12] , \A[11] , \A[10] , 
    \A[9] , \A[8] , \A[7] , \A[6] , \A[5] , \A[4] , \A[3] , \A[2] , \A[1] , \A[0] })
    , .M ({\M[31] , \M[30] , \M[29] , \M[28] , \M[27] , \M[26] , \M[25] , \M[24] , 
    \M[23] , \M[22] , \M[21] , \M[20] , \M[19] , \M[18] , \M[17] , \M[16] , \M[15] , 
    \M[14] , \M[13] , \M[12] , \M[11] , \M[10] , \M[9] , \M[8] , \M[7] , \M[6] , 
    \M[5] , \M[4] , \M[3] , \M[2] , \M[1] , \M[0] }));
datapath i_0_3 (.p_0 ({n_0_35, n_0_34, n_0_33, n_0_32, n_0_31, n_0_30, n_0_29, n_0_28, 
    n_0_27, n_0_26, n_0_25, n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, 
    n_0_17, n_0_16, n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, 
    n_0_7, n_0_6, n_0_5, n_0_4}), .A ({\A[31] , uc_0, \A[29] , \A[28] , \A[27] , 
    \A[26] , \A[25] , \A[24] , \A[23] , \A[22] , \A[21] , \A[20] , \A[19] , \A[18] , 
    \A[17] , \A[16] , \A[15] , \A[14] , \A[13] , \A[12] , \A[11] , \A[10] , \A[9] , 
    \A[8] , \A[7] , \A[6] , \A[5] , \A[4] , \A[3] , \A[2] , \A[1] , \A[0] }), .M ({
    \M[31] , \M[30] , \M[29] , \M[28] , \M[27] , \M[26] , \M[25] , \M[24] , \M[23] , 
    \M[22] , \M[21] , \M[20] , \M[19] , \M[18] , \M[17] , \M[16] , \M[15] , \M[14] , 
    \M[13] , \M[12] , \M[11] , \M[10] , \M[9] , \M[8] , \M[7] , \M[6] , \M[5] , \M[4] , 
    \M[3] , \M[2] , \M[1] , \M[0] }));
DFF_X1 \P_reg[0]  (.Q (P[0]), .CK (CTS_n105), .D (\Q[0] ));
DFF_X1 \P_reg[1]  (.Q (P[1]), .CK (CTS_n105), .D (\Q[1] ));
DFF_X1 \P_reg[2]  (.Q (P[2]), .CK (CTS_n105), .D (\Q[2] ));
DFF_X1 \P_reg[3]  (.Q (P[3]), .CK (CTS_n105), .D (\Q[3] ));
DFF_X1 \P_reg[4]  (.Q (P[4]), .CK (CTS_n105), .D (\Q[4] ));
DFF_X1 \P_reg[5]  (.Q (P[5]), .CK (CTS_n105), .D (\Q[5] ));
DFF_X1 \P_reg[6]  (.Q (P[6]), .CK (CTS_n105), .D (\Q[6] ));
DFF_X1 \P_reg[7]  (.Q (P[7]), .CK (CTS_n105), .D (\Q[7] ));
DFF_X1 \P_reg[8]  (.Q (P[8]), .CK (CTS_n105), .D (\Q[8] ));
DFF_X1 \P_reg[9]  (.Q (P[9]), .CK (CTS_n105), .D (\Q[9] ));
DFF_X1 \P_reg[10]  (.Q (P[10]), .CK (CTS_n105), .D (\Q[10] ));
DFF_X1 \P_reg[11]  (.Q (P[11]), .CK (CTS_n105), .D (\Q[11] ));
DFF_X1 \P_reg[12]  (.Q (P[12]), .CK (CTS_n105), .D (\Q[12] ));
DFF_X1 \P_reg[13]  (.Q (P[13]), .CK (CTS_n105), .D (\Q[13] ));
DFF_X1 \P_reg[14]  (.Q (P[14]), .CK (CTS_n105), .D (\Q[14] ));
DFF_X1 \P_reg[15]  (.Q (P[15]), .CK (CTS_n105), .D (\Q[15] ));
DFF_X1 \P_reg[16]  (.Q (P[16]), .CK (CTS_n105), .D (\Q[16] ));
DFF_X1 \P_reg[17]  (.Q (P[17]), .CK (CTS_n105), .D (\Q[17] ));
DFF_X1 \P_reg[18]  (.Q (P[18]), .CK (CTS_n105), .D (\Q[18] ));
DFF_X1 \P_reg[19]  (.Q (P[19]), .CK (CTS_n105), .D (\Q[19] ));
DFF_X1 \P_reg[20]  (.Q (P[20]), .CK (CTS_n105), .D (\Q[20] ));
DFF_X1 \P_reg[21]  (.Q (P[21]), .CK (CTS_n105), .D (\Q[21] ));
DFF_X1 \P_reg[22]  (.Q (P[22]), .CK (CTS_n105), .D (\Q[22] ));
DFF_X1 \P_reg[23]  (.Q (P[23]), .CK (CTS_n105), .D (\Q[23] ));
DFF_X1 \P_reg[24]  (.Q (P[24]), .CK (CTS_n105), .D (\Q[24] ));
DFF_X1 \P_reg[25]  (.Q (P[25]), .CK (CTS_n105), .D (\Q[25] ));
DFF_X1 \P_reg[26]  (.Q (P[26]), .CK (CTS_n105), .D (\Q[26] ));
DFF_X1 \P_reg[27]  (.Q (P[27]), .CK (CTS_n105), .D (\Q[27] ));
DFF_X1 \P_reg[28]  (.Q (P[28]), .CK (CTS_n105), .D (\Q[28] ));
DFF_X1 \P_reg[29]  (.Q (P[29]), .CK (CTS_n105), .D (\Q[29] ));
DFF_X1 \P_reg[30]  (.Q (P[30]), .CK (CTS_n105), .D (\Q[30] ));
DFF_X1 \P_reg[31]  (.Q (P[31]), .CK (CTS_n105), .D (\Q[31] ));
DFF_X1 \P_reg[32]  (.Q (P[32]), .CK (CTS_n105), .D (\A[0] ));
DFF_X1 \P_reg[33]  (.Q (P[33]), .CK (CTS_n105), .D (\A[1] ));
DFF_X1 \P_reg[34]  (.Q (P[34]), .CK (CTS_n105), .D (\A[2] ));
DFF_X1 \P_reg[35]  (.Q (P[35]), .CK (CTS_n105), .D (\A[3] ));
DFF_X1 \P_reg[36]  (.Q (P[36]), .CK (CTS_n105), .D (\A[4] ));
DFF_X1 \P_reg[37]  (.Q (P[37]), .CK (CTS_n105), .D (\A[5] ));
DFF_X1 \P_reg[38]  (.Q (P[38]), .CK (CTS_n105), .D (\A[6] ));
DFF_X1 \P_reg[39]  (.Q (P[39]), .CK (CTS_n105), .D (\A[7] ));
DFF_X1 \P_reg[40]  (.Q (P[40]), .CK (CTS_n105), .D (\A[8] ));
DFF_X1 \P_reg[41]  (.Q (P[41]), .CK (CTS_n105), .D (\A[9] ));
DFF_X1 \P_reg[42]  (.Q (P[42]), .CK (CTS_n105), .D (\A[10] ));
DFF_X1 \P_reg[43]  (.Q (P[43]), .CK (CTS_n105), .D (\A[11] ));
DFF_X1 \P_reg[44]  (.Q (P[44]), .CK (CTS_n105), .D (\A[12] ));
DFF_X1 \P_reg[45]  (.Q (P[45]), .CK (CTS_n105), .D (\A[13] ));
DFF_X1 \P_reg[46]  (.Q (P[46]), .CK (CTS_n105), .D (\A[14] ));
DFF_X1 \P_reg[47]  (.Q (P[47]), .CK (CTS_n105), .D (\A[15] ));
DFF_X1 \P_reg[48]  (.Q (P[48]), .CK (CTS_n105), .D (\A[16] ));
DFF_X1 \P_reg[49]  (.Q (P[49]), .CK (CTS_n105), .D (\A[17] ));
DFF_X1 \P_reg[50]  (.Q (P[50]), .CK (CTS_n105), .D (\A[18] ));
DFF_X1 \P_reg[51]  (.Q (P[51]), .CK (CTS_n105), .D (\A[19] ));
DFF_X1 \P_reg[52]  (.Q (P[52]), .CK (CTS_n105), .D (\A[20] ));
DFF_X1 \P_reg[53]  (.Q (P[53]), .CK (CTS_n105), .D (\A[21] ));
DFF_X1 \P_reg[54]  (.Q (P[54]), .CK (CTS_n105), .D (\A[22] ));
DFF_X1 \P_reg[55]  (.Q (P[55]), .CK (CTS_n105), .D (\A[23] ));
DFF_X1 \P_reg[56]  (.Q (P[56]), .CK (CTS_n105), .D (\A[24] ));
DFF_X1 \P_reg[57]  (.Q (P[57]), .CK (CTS_n105), .D (\A[25] ));
DFF_X1 \P_reg[58]  (.Q (P[58]), .CK (CTS_n105), .D (\A[26] ));
DFF_X1 \P_reg[59]  (.Q (P[59]), .CK (CTS_n105), .D (\A[27] ));
DFF_X1 \P_reg[60]  (.Q (P[60]), .CK (CTS_n105), .D (\A[28] ));
DFF_X1 \P_reg[61]  (.Q (P[61]), .CK (CTS_n105), .D (\A[29] ));
DFF_X1 \P_reg[63]  (.Q (P[62]), .CK (CTS_n105), .D (\A[31] ));
CLKGATETST_X8 clk_gate_P_reg (.GCK (CTS_n106), .CK (clk), .E (n_0_104), .SE (1'b0 ));
CLKBUF_X2 drc_ipo_c6 (.Z (drc_ipo_n6), .A (n_0_0_33));
CLKBUF_X2 drc_ipo_c5 (.Z (drc_ipo_n5), .A (n_0_0_34));
CLKBUF_X3 CTS_L3_c11 (.Z (CTS_n8), .A (CTS_n56));
CLKBUF_X3 CTS_L3_c12 (.Z (CTS_n9), .A (CTS_n56));
CLKBUF_X3 CTS_L2_c73 (.Z (CTS_n105), .A (CTS_n106));
CLKBUF_X1 CTS_L1_c148 (.Z (CTS_n214), .A (clk));
CLKBUF_X1 CTS_L2_c129 (.Z (CTS_n178), .A (CTS_n214));
CLKBUF_X2 CTS_L1_c142 (.Z (CTS_n193), .A (clk));
CLKBUF_X1 CLOCK_slh__c151 (.Z (CLOCK_slh_n243), .A (m[17]));
CLKBUF_X1 CLOCK_slh__c153 (.Z (CLOCK_slh_n248), .A (m[18]));
CLKBUF_X1 CLOCK_slh__c155 (.Z (CLOCK_slh_n253), .A (m[20]));
CLKBUF_X1 CLOCK_slh__c157 (.Z (CLOCK_slh_n258), .A (m[21]));
CLKBUF_X1 CLOCK_slh__c159 (.Z (CLOCK_slh_n263), .A (m[12]));
CLKBUF_X1 CLOCK_slh__c161 (.Z (CLOCK_slh_n268), .A (m[16]));
CLKBUF_X1 CLOCK_slh__c163 (.Z (CLOCK_slh_n273), .A (m[22]));
CLKBUF_X1 CLOCK_slh__c165 (.Z (CLOCK_slh_n278), .A (m[23]));
CLKBUF_X1 CLOCK_slh__c167 (.Z (CLOCK_slh_n283), .A (m[15]));
CLKBUF_X1 CLOCK_slh__c169 (.Z (CLOCK_slh_n288), .A (m[7]));
CLKBUF_X1 CLOCK_slh__c171 (.Z (CLOCK_slh_n293), .A (m[31]));
CLKBUF_X1 CLOCK_slh__c173 (.Z (CLOCK_slh_n298), .A (m[19]));
CLKBUF_X1 CLOCK_slh__c175 (.Z (CLOCK_slh_n303), .A (m[8]));
CLKBUF_X1 CLOCK_slh__c177 (.Z (CLOCK_slh_n308), .A (m[3]));
CLKBUF_X1 CLOCK_slh__c179 (.Z (CLOCK_slh_n313), .A (m[5]));
CLKBUF_X1 CLOCK_slh__c181 (.Z (CLOCK_slh_n318), .A (m[10]));
CLKBUF_X1 CLOCK_slh__c183 (.Z (CLOCK_slh_n323), .A (m[11]));
CLKBUF_X1 CLOCK_slh__c185 (.Z (CLOCK_slh_n328), .A (m[13]));
CLKBUF_X1 CLOCK_slh__c187 (.Z (CLOCK_slh_n333), .A (m[14]));
CLKBUF_X1 CLOCK_slh__c189 (.Z (CLOCK_slh_n338), .A (m[4]));
CLKBUF_X1 CLOCK_slh__c191 (.Z (CLOCK_slh_n343), .A (m[6]));
CLKBUF_X1 CLOCK_slh__c193 (.Z (CLOCK_slh_n348), .A (m[9]));
CLKBUF_X1 CLOCK_slh__c195 (.Z (CLOCK_slh_n353), .A (m[2]));
CLKBUF_X1 CLOCK_slh__c197 (.Z (CLOCK_slh_n358), .A (m[1]));
CLKBUF_X1 CLOCK_slh__c199 (.Z (CLOCK_slh_n363), .A (m[0]));
CLKBUF_X1 CLOCK_slh__c201 (.Z (CLOCK_slh_n368), .A (m[26]));
CLKBUF_X1 CLOCK_slh__c203 (.Z (CLOCK_slh_n373), .A (m[30]));
CLKBUF_X1 CLOCK_slh__c205 (.Z (CLOCK_slh_n378), .A (m[24]));
CLKBUF_X1 CLOCK_slh__c207 (.Z (CLOCK_slh_n383), .A (m[28]));
CLKBUF_X1 CLOCK_slh__c209 (.Z (CLOCK_slh_n388), .A (m[25]));
CLKBUF_X1 CLOCK_slh__c211 (.Z (CLOCK_slh_n393), .A (m[29]));
CLKBUF_X1 CLOCK_slh__c213 (.Z (CLOCK_slh_n398), .A (m[27]));

endmodule //Booth


